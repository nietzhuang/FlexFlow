module Bank(
  input         clock,
  input         reset,
  input  [15:0] io_BankIO_DataIn,
  input  [9:0]  io_BankIO_DataAddr,
  input         io_BankIO_ReadWrite,
  input         io_BankIO_Enable,
  output [15:0] io_BankIO_DataOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] buffer_0; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_2; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_3; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_4; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_5; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_6; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_7; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_8; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_9; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_10; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_11; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_12; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_13; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_14; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_15; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_16; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_17; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_18; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_19; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_20; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_21; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_22; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_23; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_24; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_25; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_26; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_27; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_28; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_29; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_30; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_31; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_32; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_33; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_34; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_35; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_36; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_37; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_38; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_39; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_40; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_41; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_42; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_43; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_44; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_45; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_46; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_47; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_48; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_49; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_50; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_51; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_52; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_53; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_54; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_55; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_56; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_57; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_58; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_59; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_60; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_61; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_62; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_63; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_64; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_65; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_66; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_67; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_68; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_69; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_70; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_71; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_72; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_73; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_74; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_75; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_76; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_77; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_78; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_79; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_80; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_81; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_82; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_83; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_84; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_85; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_86; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_87; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_88; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_89; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_90; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_91; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_92; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_93; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_94; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_95; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_96; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_97; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_98; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_99; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_100; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_101; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_102; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_103; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_104; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_105; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_106; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_107; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_108; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_109; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_110; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_111; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_112; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_113; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_114; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_115; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_116; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_117; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_118; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_119; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_120; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_121; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_122; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_123; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_124; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_125; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_126; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_127; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_128; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_129; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_130; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_131; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_132; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_133; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_134; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_135; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_136; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_137; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_138; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_139; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_140; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_141; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_142; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_143; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_144; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_145; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_146; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_147; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_148; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_149; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_150; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_151; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_152; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_153; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_154; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_155; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_156; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_157; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_158; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_159; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_160; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_161; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_162; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_163; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_164; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_165; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_166; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_167; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_168; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_169; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_170; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_171; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_172; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_173; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_174; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_175; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_176; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_177; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_178; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_179; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_180; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_181; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_182; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_183; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_184; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_185; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_186; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_187; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_188; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_189; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_190; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_191; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_192; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_193; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_194; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_195; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_196; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_197; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_198; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_199; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_200; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_201; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_202; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_203; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_204; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_205; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_206; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_207; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_208; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_209; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_210; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_211; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_212; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_213; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_214; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_215; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_216; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_217; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_218; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_219; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_220; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_221; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_222; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_223; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_224; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_225; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_226; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_227; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_228; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_229; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_230; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_231; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_232; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_233; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_234; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_235; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_236; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_237; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_238; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_239; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_240; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_241; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_242; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_243; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_244; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_245; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_246; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_247; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_248; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_249; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_250; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_251; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_252; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_253; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_254; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_255; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_256; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_257; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_258; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_259; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_260; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_261; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_262; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_263; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_264; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_265; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_266; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_267; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_268; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_269; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_270; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_271; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_272; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_273; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_274; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_275; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_276; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_277; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_278; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_279; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_280; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_281; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_282; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_283; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_284; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_285; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_286; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_287; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_288; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_289; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_290; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_291; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_292; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_293; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_294; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_295; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_296; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_297; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_298; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_299; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_300; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_301; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_302; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_303; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_304; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_305; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_306; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_307; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_308; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_309; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_310; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_311; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_312; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_313; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_314; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_315; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_316; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_317; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_318; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_319; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_320; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_321; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_322; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_323; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_324; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_325; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_326; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_327; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_328; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_329; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_330; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_331; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_332; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_333; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_334; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_335; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_336; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_337; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_338; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_339; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_340; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_341; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_342; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_343; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_344; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_345; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_346; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_347; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_348; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_349; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_350; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_351; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_352; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_353; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_354; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_355; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_356; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_357; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_358; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_359; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_360; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_361; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_362; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_363; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_364; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_365; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_366; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_367; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_368; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_369; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_370; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_371; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_372; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_373; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_374; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_375; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_376; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_377; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_378; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_379; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_380; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_381; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_382; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_383; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_384; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_385; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_386; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_387; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_388; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_389; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_390; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_391; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_392; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_393; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_394; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_395; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_396; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_397; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_398; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_399; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_400; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_401; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_402; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_403; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_404; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_405; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_406; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_407; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_408; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_409; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_410; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_411; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_412; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_413; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_414; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_415; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_416; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_417; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_418; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_419; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_420; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_421; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_422; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_423; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_424; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_425; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_426; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_427; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_428; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_429; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_430; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_431; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_432; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_433; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_434; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_435; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_436; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_437; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_438; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_439; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_440; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_441; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_442; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_443; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_444; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_445; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_446; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_447; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_448; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_449; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_450; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_451; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_452; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_453; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_454; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_455; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_456; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_457; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_458; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_459; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_460; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_461; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_462; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_463; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_464; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_465; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_466; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_467; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_468; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_469; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_470; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_471; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_472; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_473; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_474; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_475; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_476; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_477; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_478; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_479; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_480; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_481; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_482; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_483; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_484; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_485; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_486; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_487; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_488; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_489; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_490; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_491; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_492; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_493; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_494; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_495; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_496; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_497; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_498; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_499; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_500; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_501; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_502; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_503; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_504; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_505; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_506; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_507; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_508; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_509; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_510; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_511; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_512; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_513; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_514; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_515; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_516; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_517; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_518; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_519; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_520; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_521; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_522; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_523; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_524; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_525; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_526; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_527; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_528; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_529; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_530; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_531; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_532; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_533; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_534; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_535; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_536; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_537; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_538; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_539; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_540; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_541; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_542; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_543; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_544; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_545; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_546; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_547; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_548; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_549; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_550; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_551; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_552; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_553; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_554; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_555; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_556; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_557; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_558; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_559; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_560; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_561; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_562; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_563; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_564; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_565; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_566; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_567; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_568; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_569; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_570; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_571; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_572; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_573; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_574; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_575; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_576; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_577; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_578; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_579; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_580; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_581; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_582; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_583; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_584; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_585; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_586; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_587; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_588; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_589; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_590; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_591; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_592; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_593; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_594; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_595; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_596; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_597; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_598; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_599; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_600; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_601; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_602; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_603; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_604; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_605; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_606; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_607; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_608; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_609; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_610; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_611; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_612; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_613; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_614; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_615; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_616; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_617; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_618; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_619; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_620; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_621; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_622; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_623; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_624; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_625; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_626; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_627; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_628; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_629; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_630; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_631; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_632; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_633; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_634; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_635; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_636; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_637; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_638; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_639; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_640; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_641; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_642; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_643; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_644; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_645; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_646; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_647; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_648; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_649; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_650; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_651; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_652; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_653; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_654; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_655; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_656; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_657; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_658; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_659; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_660; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_661; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_662; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_663; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_664; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_665; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_666; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_667; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_668; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_669; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_670; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_671; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_672; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_673; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_674; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_675; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_676; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_677; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_678; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_679; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_680; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_681; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_682; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_683; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_684; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_685; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_686; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_687; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_688; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_689; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_690; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_691; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_692; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_693; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_694; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_695; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_696; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_697; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_698; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_699; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_700; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_701; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_702; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_703; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_704; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_705; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_706; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_707; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_708; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_709; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_710; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_711; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_712; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_713; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_714; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_715; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_716; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_717; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_718; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_719; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_720; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_721; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_722; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_723; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_724; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_725; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_726; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_727; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_728; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_729; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_730; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_731; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_732; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_733; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_734; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_735; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_736; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_737; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_738; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_739; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_740; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_741; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_742; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_743; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_744; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_745; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_746; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_747; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_748; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_749; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_750; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_751; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_752; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_753; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_754; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_755; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_756; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_757; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_758; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_759; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_760; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_761; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_762; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_763; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_764; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_765; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_766; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_767; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_768; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_769; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_770; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_771; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_772; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_773; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_774; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_775; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_776; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_777; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_778; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_779; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_780; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_781; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_782; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_783; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_784; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_785; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_786; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_787; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_788; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_789; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_790; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_791; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_792; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_793; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_794; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_795; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_796; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_797; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_798; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_799; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_800; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_801; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_802; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_803; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_804; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_805; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_806; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_807; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_808; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_809; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_810; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_811; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_812; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_813; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_814; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_815; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_816; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_817; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_818; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_819; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_820; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_821; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_822; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_823; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_824; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_825; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_826; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_827; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_828; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_829; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_830; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_831; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_832; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_833; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_834; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_835; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_836; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_837; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_838; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_839; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_840; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_841; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_842; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_843; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_844; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_845; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_846; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_847; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_848; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_849; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_850; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_851; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_852; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_853; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_854; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_855; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_856; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_857; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_858; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_859; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_860; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_861; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_862; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_863; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_864; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_865; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_866; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_867; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_868; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_869; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_870; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_871; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_872; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_873; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_874; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_875; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_876; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_877; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_878; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_879; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_880; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_881; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_882; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_883; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_884; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_885; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_886; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_887; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_888; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_889; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_890; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_891; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_892; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_893; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_894; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_895; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_896; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_897; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_898; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_899; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_900; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_901; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_902; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_903; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_904; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_905; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_906; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_907; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_908; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_909; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_910; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_911; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_912; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_913; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_914; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_915; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_916; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_917; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_918; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_919; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_920; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_921; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_922; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_923; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_924; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_925; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_926; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_927; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_928; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_929; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_930; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_931; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_932; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_933; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_934; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_935; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_936; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_937; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_938; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_939; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_940; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_941; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_942; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_943; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_944; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_945; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_946; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_947; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_948; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_949; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_950; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_951; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_952; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_953; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_954; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_955; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_956; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_957; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_958; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_959; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_960; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_961; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_962; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_963; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_964; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_965; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_966; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_967; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_968; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_969; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_970; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_971; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_972; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_973; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_974; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_975; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_976; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_977; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_978; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_979; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_980; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_981; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_982; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_983; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_984; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_985; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_986; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_987; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_988; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_989; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_990; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_991; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_992; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_993; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_994; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_995; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_996; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_997; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_998; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_999; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1000; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1001; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1002; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1003; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1004; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1005; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1006; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1007; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1008; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1009; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1010; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1011; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1012; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1013; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1014; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1015; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1016; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1017; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1018; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1019; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1020; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1021; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1022; // @[OuterBuffer.scala 20:24]
  reg [15:0] buffer_1023; // @[OuterBuffer.scala 20:24]
  wire [15:0] _GEN_1025 = 10'h1 == io_BankIO_DataAddr ? buffer_1 : buffer_0; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1026 = 10'h2 == io_BankIO_DataAddr ? buffer_2 : _GEN_1025; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1027 = 10'h3 == io_BankIO_DataAddr ? buffer_3 : _GEN_1026; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1028 = 10'h4 == io_BankIO_DataAddr ? buffer_4 : _GEN_1027; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1029 = 10'h5 == io_BankIO_DataAddr ? buffer_5 : _GEN_1028; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1030 = 10'h6 == io_BankIO_DataAddr ? buffer_6 : _GEN_1029; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1031 = 10'h7 == io_BankIO_DataAddr ? buffer_7 : _GEN_1030; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1032 = 10'h8 == io_BankIO_DataAddr ? buffer_8 : _GEN_1031; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1033 = 10'h9 == io_BankIO_DataAddr ? buffer_9 : _GEN_1032; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1034 = 10'ha == io_BankIO_DataAddr ? buffer_10 : _GEN_1033; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1035 = 10'hb == io_BankIO_DataAddr ? buffer_11 : _GEN_1034; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1036 = 10'hc == io_BankIO_DataAddr ? buffer_12 : _GEN_1035; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1037 = 10'hd == io_BankIO_DataAddr ? buffer_13 : _GEN_1036; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1038 = 10'he == io_BankIO_DataAddr ? buffer_14 : _GEN_1037; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1039 = 10'hf == io_BankIO_DataAddr ? buffer_15 : _GEN_1038; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1040 = 10'h10 == io_BankIO_DataAddr ? buffer_16 : _GEN_1039; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1041 = 10'h11 == io_BankIO_DataAddr ? buffer_17 : _GEN_1040; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1042 = 10'h12 == io_BankIO_DataAddr ? buffer_18 : _GEN_1041; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1043 = 10'h13 == io_BankIO_DataAddr ? buffer_19 : _GEN_1042; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1044 = 10'h14 == io_BankIO_DataAddr ? buffer_20 : _GEN_1043; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1045 = 10'h15 == io_BankIO_DataAddr ? buffer_21 : _GEN_1044; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1046 = 10'h16 == io_BankIO_DataAddr ? buffer_22 : _GEN_1045; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1047 = 10'h17 == io_BankIO_DataAddr ? buffer_23 : _GEN_1046; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1048 = 10'h18 == io_BankIO_DataAddr ? buffer_24 : _GEN_1047; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1049 = 10'h19 == io_BankIO_DataAddr ? buffer_25 : _GEN_1048; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1050 = 10'h1a == io_BankIO_DataAddr ? buffer_26 : _GEN_1049; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1051 = 10'h1b == io_BankIO_DataAddr ? buffer_27 : _GEN_1050; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1052 = 10'h1c == io_BankIO_DataAddr ? buffer_28 : _GEN_1051; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1053 = 10'h1d == io_BankIO_DataAddr ? buffer_29 : _GEN_1052; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1054 = 10'h1e == io_BankIO_DataAddr ? buffer_30 : _GEN_1053; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1055 = 10'h1f == io_BankIO_DataAddr ? buffer_31 : _GEN_1054; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1056 = 10'h20 == io_BankIO_DataAddr ? buffer_32 : _GEN_1055; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1057 = 10'h21 == io_BankIO_DataAddr ? buffer_33 : _GEN_1056; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1058 = 10'h22 == io_BankIO_DataAddr ? buffer_34 : _GEN_1057; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1059 = 10'h23 == io_BankIO_DataAddr ? buffer_35 : _GEN_1058; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1060 = 10'h24 == io_BankIO_DataAddr ? buffer_36 : _GEN_1059; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1061 = 10'h25 == io_BankIO_DataAddr ? buffer_37 : _GEN_1060; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1062 = 10'h26 == io_BankIO_DataAddr ? buffer_38 : _GEN_1061; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1063 = 10'h27 == io_BankIO_DataAddr ? buffer_39 : _GEN_1062; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1064 = 10'h28 == io_BankIO_DataAddr ? buffer_40 : _GEN_1063; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1065 = 10'h29 == io_BankIO_DataAddr ? buffer_41 : _GEN_1064; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1066 = 10'h2a == io_BankIO_DataAddr ? buffer_42 : _GEN_1065; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1067 = 10'h2b == io_BankIO_DataAddr ? buffer_43 : _GEN_1066; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1068 = 10'h2c == io_BankIO_DataAddr ? buffer_44 : _GEN_1067; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1069 = 10'h2d == io_BankIO_DataAddr ? buffer_45 : _GEN_1068; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1070 = 10'h2e == io_BankIO_DataAddr ? buffer_46 : _GEN_1069; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1071 = 10'h2f == io_BankIO_DataAddr ? buffer_47 : _GEN_1070; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1072 = 10'h30 == io_BankIO_DataAddr ? buffer_48 : _GEN_1071; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1073 = 10'h31 == io_BankIO_DataAddr ? buffer_49 : _GEN_1072; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1074 = 10'h32 == io_BankIO_DataAddr ? buffer_50 : _GEN_1073; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1075 = 10'h33 == io_BankIO_DataAddr ? buffer_51 : _GEN_1074; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1076 = 10'h34 == io_BankIO_DataAddr ? buffer_52 : _GEN_1075; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1077 = 10'h35 == io_BankIO_DataAddr ? buffer_53 : _GEN_1076; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1078 = 10'h36 == io_BankIO_DataAddr ? buffer_54 : _GEN_1077; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1079 = 10'h37 == io_BankIO_DataAddr ? buffer_55 : _GEN_1078; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1080 = 10'h38 == io_BankIO_DataAddr ? buffer_56 : _GEN_1079; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1081 = 10'h39 == io_BankIO_DataAddr ? buffer_57 : _GEN_1080; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1082 = 10'h3a == io_BankIO_DataAddr ? buffer_58 : _GEN_1081; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1083 = 10'h3b == io_BankIO_DataAddr ? buffer_59 : _GEN_1082; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1084 = 10'h3c == io_BankIO_DataAddr ? buffer_60 : _GEN_1083; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1085 = 10'h3d == io_BankIO_DataAddr ? buffer_61 : _GEN_1084; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1086 = 10'h3e == io_BankIO_DataAddr ? buffer_62 : _GEN_1085; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1087 = 10'h3f == io_BankIO_DataAddr ? buffer_63 : _GEN_1086; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1088 = 10'h40 == io_BankIO_DataAddr ? buffer_64 : _GEN_1087; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1089 = 10'h41 == io_BankIO_DataAddr ? buffer_65 : _GEN_1088; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1090 = 10'h42 == io_BankIO_DataAddr ? buffer_66 : _GEN_1089; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1091 = 10'h43 == io_BankIO_DataAddr ? buffer_67 : _GEN_1090; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1092 = 10'h44 == io_BankIO_DataAddr ? buffer_68 : _GEN_1091; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1093 = 10'h45 == io_BankIO_DataAddr ? buffer_69 : _GEN_1092; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1094 = 10'h46 == io_BankIO_DataAddr ? buffer_70 : _GEN_1093; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1095 = 10'h47 == io_BankIO_DataAddr ? buffer_71 : _GEN_1094; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1096 = 10'h48 == io_BankIO_DataAddr ? buffer_72 : _GEN_1095; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1097 = 10'h49 == io_BankIO_DataAddr ? buffer_73 : _GEN_1096; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1098 = 10'h4a == io_BankIO_DataAddr ? buffer_74 : _GEN_1097; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1099 = 10'h4b == io_BankIO_DataAddr ? buffer_75 : _GEN_1098; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1100 = 10'h4c == io_BankIO_DataAddr ? buffer_76 : _GEN_1099; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1101 = 10'h4d == io_BankIO_DataAddr ? buffer_77 : _GEN_1100; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1102 = 10'h4e == io_BankIO_DataAddr ? buffer_78 : _GEN_1101; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1103 = 10'h4f == io_BankIO_DataAddr ? buffer_79 : _GEN_1102; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1104 = 10'h50 == io_BankIO_DataAddr ? buffer_80 : _GEN_1103; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1105 = 10'h51 == io_BankIO_DataAddr ? buffer_81 : _GEN_1104; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1106 = 10'h52 == io_BankIO_DataAddr ? buffer_82 : _GEN_1105; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1107 = 10'h53 == io_BankIO_DataAddr ? buffer_83 : _GEN_1106; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1108 = 10'h54 == io_BankIO_DataAddr ? buffer_84 : _GEN_1107; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1109 = 10'h55 == io_BankIO_DataAddr ? buffer_85 : _GEN_1108; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1110 = 10'h56 == io_BankIO_DataAddr ? buffer_86 : _GEN_1109; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1111 = 10'h57 == io_BankIO_DataAddr ? buffer_87 : _GEN_1110; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1112 = 10'h58 == io_BankIO_DataAddr ? buffer_88 : _GEN_1111; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1113 = 10'h59 == io_BankIO_DataAddr ? buffer_89 : _GEN_1112; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1114 = 10'h5a == io_BankIO_DataAddr ? buffer_90 : _GEN_1113; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1115 = 10'h5b == io_BankIO_DataAddr ? buffer_91 : _GEN_1114; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1116 = 10'h5c == io_BankIO_DataAddr ? buffer_92 : _GEN_1115; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1117 = 10'h5d == io_BankIO_DataAddr ? buffer_93 : _GEN_1116; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1118 = 10'h5e == io_BankIO_DataAddr ? buffer_94 : _GEN_1117; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1119 = 10'h5f == io_BankIO_DataAddr ? buffer_95 : _GEN_1118; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1120 = 10'h60 == io_BankIO_DataAddr ? buffer_96 : _GEN_1119; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1121 = 10'h61 == io_BankIO_DataAddr ? buffer_97 : _GEN_1120; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1122 = 10'h62 == io_BankIO_DataAddr ? buffer_98 : _GEN_1121; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1123 = 10'h63 == io_BankIO_DataAddr ? buffer_99 : _GEN_1122; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1124 = 10'h64 == io_BankIO_DataAddr ? buffer_100 : _GEN_1123; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1125 = 10'h65 == io_BankIO_DataAddr ? buffer_101 : _GEN_1124; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1126 = 10'h66 == io_BankIO_DataAddr ? buffer_102 : _GEN_1125; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1127 = 10'h67 == io_BankIO_DataAddr ? buffer_103 : _GEN_1126; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1128 = 10'h68 == io_BankIO_DataAddr ? buffer_104 : _GEN_1127; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1129 = 10'h69 == io_BankIO_DataAddr ? buffer_105 : _GEN_1128; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1130 = 10'h6a == io_BankIO_DataAddr ? buffer_106 : _GEN_1129; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1131 = 10'h6b == io_BankIO_DataAddr ? buffer_107 : _GEN_1130; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1132 = 10'h6c == io_BankIO_DataAddr ? buffer_108 : _GEN_1131; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1133 = 10'h6d == io_BankIO_DataAddr ? buffer_109 : _GEN_1132; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1134 = 10'h6e == io_BankIO_DataAddr ? buffer_110 : _GEN_1133; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1135 = 10'h6f == io_BankIO_DataAddr ? buffer_111 : _GEN_1134; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1136 = 10'h70 == io_BankIO_DataAddr ? buffer_112 : _GEN_1135; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1137 = 10'h71 == io_BankIO_DataAddr ? buffer_113 : _GEN_1136; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1138 = 10'h72 == io_BankIO_DataAddr ? buffer_114 : _GEN_1137; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1139 = 10'h73 == io_BankIO_DataAddr ? buffer_115 : _GEN_1138; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1140 = 10'h74 == io_BankIO_DataAddr ? buffer_116 : _GEN_1139; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1141 = 10'h75 == io_BankIO_DataAddr ? buffer_117 : _GEN_1140; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1142 = 10'h76 == io_BankIO_DataAddr ? buffer_118 : _GEN_1141; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1143 = 10'h77 == io_BankIO_DataAddr ? buffer_119 : _GEN_1142; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1144 = 10'h78 == io_BankIO_DataAddr ? buffer_120 : _GEN_1143; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1145 = 10'h79 == io_BankIO_DataAddr ? buffer_121 : _GEN_1144; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1146 = 10'h7a == io_BankIO_DataAddr ? buffer_122 : _GEN_1145; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1147 = 10'h7b == io_BankIO_DataAddr ? buffer_123 : _GEN_1146; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1148 = 10'h7c == io_BankIO_DataAddr ? buffer_124 : _GEN_1147; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1149 = 10'h7d == io_BankIO_DataAddr ? buffer_125 : _GEN_1148; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1150 = 10'h7e == io_BankIO_DataAddr ? buffer_126 : _GEN_1149; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1151 = 10'h7f == io_BankIO_DataAddr ? buffer_127 : _GEN_1150; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1152 = 10'h80 == io_BankIO_DataAddr ? buffer_128 : _GEN_1151; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1153 = 10'h81 == io_BankIO_DataAddr ? buffer_129 : _GEN_1152; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1154 = 10'h82 == io_BankIO_DataAddr ? buffer_130 : _GEN_1153; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1155 = 10'h83 == io_BankIO_DataAddr ? buffer_131 : _GEN_1154; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1156 = 10'h84 == io_BankIO_DataAddr ? buffer_132 : _GEN_1155; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1157 = 10'h85 == io_BankIO_DataAddr ? buffer_133 : _GEN_1156; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1158 = 10'h86 == io_BankIO_DataAddr ? buffer_134 : _GEN_1157; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1159 = 10'h87 == io_BankIO_DataAddr ? buffer_135 : _GEN_1158; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1160 = 10'h88 == io_BankIO_DataAddr ? buffer_136 : _GEN_1159; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1161 = 10'h89 == io_BankIO_DataAddr ? buffer_137 : _GEN_1160; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1162 = 10'h8a == io_BankIO_DataAddr ? buffer_138 : _GEN_1161; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1163 = 10'h8b == io_BankIO_DataAddr ? buffer_139 : _GEN_1162; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1164 = 10'h8c == io_BankIO_DataAddr ? buffer_140 : _GEN_1163; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1165 = 10'h8d == io_BankIO_DataAddr ? buffer_141 : _GEN_1164; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1166 = 10'h8e == io_BankIO_DataAddr ? buffer_142 : _GEN_1165; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1167 = 10'h8f == io_BankIO_DataAddr ? buffer_143 : _GEN_1166; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1168 = 10'h90 == io_BankIO_DataAddr ? buffer_144 : _GEN_1167; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1169 = 10'h91 == io_BankIO_DataAddr ? buffer_145 : _GEN_1168; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1170 = 10'h92 == io_BankIO_DataAddr ? buffer_146 : _GEN_1169; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1171 = 10'h93 == io_BankIO_DataAddr ? buffer_147 : _GEN_1170; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1172 = 10'h94 == io_BankIO_DataAddr ? buffer_148 : _GEN_1171; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1173 = 10'h95 == io_BankIO_DataAddr ? buffer_149 : _GEN_1172; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1174 = 10'h96 == io_BankIO_DataAddr ? buffer_150 : _GEN_1173; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1175 = 10'h97 == io_BankIO_DataAddr ? buffer_151 : _GEN_1174; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1176 = 10'h98 == io_BankIO_DataAddr ? buffer_152 : _GEN_1175; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1177 = 10'h99 == io_BankIO_DataAddr ? buffer_153 : _GEN_1176; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1178 = 10'h9a == io_BankIO_DataAddr ? buffer_154 : _GEN_1177; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1179 = 10'h9b == io_BankIO_DataAddr ? buffer_155 : _GEN_1178; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1180 = 10'h9c == io_BankIO_DataAddr ? buffer_156 : _GEN_1179; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1181 = 10'h9d == io_BankIO_DataAddr ? buffer_157 : _GEN_1180; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1182 = 10'h9e == io_BankIO_DataAddr ? buffer_158 : _GEN_1181; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1183 = 10'h9f == io_BankIO_DataAddr ? buffer_159 : _GEN_1182; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1184 = 10'ha0 == io_BankIO_DataAddr ? buffer_160 : _GEN_1183; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1185 = 10'ha1 == io_BankIO_DataAddr ? buffer_161 : _GEN_1184; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1186 = 10'ha2 == io_BankIO_DataAddr ? buffer_162 : _GEN_1185; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1187 = 10'ha3 == io_BankIO_DataAddr ? buffer_163 : _GEN_1186; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1188 = 10'ha4 == io_BankIO_DataAddr ? buffer_164 : _GEN_1187; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1189 = 10'ha5 == io_BankIO_DataAddr ? buffer_165 : _GEN_1188; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1190 = 10'ha6 == io_BankIO_DataAddr ? buffer_166 : _GEN_1189; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1191 = 10'ha7 == io_BankIO_DataAddr ? buffer_167 : _GEN_1190; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1192 = 10'ha8 == io_BankIO_DataAddr ? buffer_168 : _GEN_1191; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1193 = 10'ha9 == io_BankIO_DataAddr ? buffer_169 : _GEN_1192; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1194 = 10'haa == io_BankIO_DataAddr ? buffer_170 : _GEN_1193; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1195 = 10'hab == io_BankIO_DataAddr ? buffer_171 : _GEN_1194; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1196 = 10'hac == io_BankIO_DataAddr ? buffer_172 : _GEN_1195; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1197 = 10'had == io_BankIO_DataAddr ? buffer_173 : _GEN_1196; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1198 = 10'hae == io_BankIO_DataAddr ? buffer_174 : _GEN_1197; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1199 = 10'haf == io_BankIO_DataAddr ? buffer_175 : _GEN_1198; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1200 = 10'hb0 == io_BankIO_DataAddr ? buffer_176 : _GEN_1199; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1201 = 10'hb1 == io_BankIO_DataAddr ? buffer_177 : _GEN_1200; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1202 = 10'hb2 == io_BankIO_DataAddr ? buffer_178 : _GEN_1201; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1203 = 10'hb3 == io_BankIO_DataAddr ? buffer_179 : _GEN_1202; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1204 = 10'hb4 == io_BankIO_DataAddr ? buffer_180 : _GEN_1203; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1205 = 10'hb5 == io_BankIO_DataAddr ? buffer_181 : _GEN_1204; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1206 = 10'hb6 == io_BankIO_DataAddr ? buffer_182 : _GEN_1205; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1207 = 10'hb7 == io_BankIO_DataAddr ? buffer_183 : _GEN_1206; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1208 = 10'hb8 == io_BankIO_DataAddr ? buffer_184 : _GEN_1207; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1209 = 10'hb9 == io_BankIO_DataAddr ? buffer_185 : _GEN_1208; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1210 = 10'hba == io_BankIO_DataAddr ? buffer_186 : _GEN_1209; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1211 = 10'hbb == io_BankIO_DataAddr ? buffer_187 : _GEN_1210; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1212 = 10'hbc == io_BankIO_DataAddr ? buffer_188 : _GEN_1211; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1213 = 10'hbd == io_BankIO_DataAddr ? buffer_189 : _GEN_1212; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1214 = 10'hbe == io_BankIO_DataAddr ? buffer_190 : _GEN_1213; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1215 = 10'hbf == io_BankIO_DataAddr ? buffer_191 : _GEN_1214; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1216 = 10'hc0 == io_BankIO_DataAddr ? buffer_192 : _GEN_1215; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1217 = 10'hc1 == io_BankIO_DataAddr ? buffer_193 : _GEN_1216; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1218 = 10'hc2 == io_BankIO_DataAddr ? buffer_194 : _GEN_1217; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1219 = 10'hc3 == io_BankIO_DataAddr ? buffer_195 : _GEN_1218; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1220 = 10'hc4 == io_BankIO_DataAddr ? buffer_196 : _GEN_1219; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1221 = 10'hc5 == io_BankIO_DataAddr ? buffer_197 : _GEN_1220; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1222 = 10'hc6 == io_BankIO_DataAddr ? buffer_198 : _GEN_1221; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1223 = 10'hc7 == io_BankIO_DataAddr ? buffer_199 : _GEN_1222; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1224 = 10'hc8 == io_BankIO_DataAddr ? buffer_200 : _GEN_1223; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1225 = 10'hc9 == io_BankIO_DataAddr ? buffer_201 : _GEN_1224; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1226 = 10'hca == io_BankIO_DataAddr ? buffer_202 : _GEN_1225; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1227 = 10'hcb == io_BankIO_DataAddr ? buffer_203 : _GEN_1226; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1228 = 10'hcc == io_BankIO_DataAddr ? buffer_204 : _GEN_1227; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1229 = 10'hcd == io_BankIO_DataAddr ? buffer_205 : _GEN_1228; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1230 = 10'hce == io_BankIO_DataAddr ? buffer_206 : _GEN_1229; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1231 = 10'hcf == io_BankIO_DataAddr ? buffer_207 : _GEN_1230; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1232 = 10'hd0 == io_BankIO_DataAddr ? buffer_208 : _GEN_1231; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1233 = 10'hd1 == io_BankIO_DataAddr ? buffer_209 : _GEN_1232; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1234 = 10'hd2 == io_BankIO_DataAddr ? buffer_210 : _GEN_1233; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1235 = 10'hd3 == io_BankIO_DataAddr ? buffer_211 : _GEN_1234; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1236 = 10'hd4 == io_BankIO_DataAddr ? buffer_212 : _GEN_1235; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1237 = 10'hd5 == io_BankIO_DataAddr ? buffer_213 : _GEN_1236; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1238 = 10'hd6 == io_BankIO_DataAddr ? buffer_214 : _GEN_1237; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1239 = 10'hd7 == io_BankIO_DataAddr ? buffer_215 : _GEN_1238; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1240 = 10'hd8 == io_BankIO_DataAddr ? buffer_216 : _GEN_1239; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1241 = 10'hd9 == io_BankIO_DataAddr ? buffer_217 : _GEN_1240; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1242 = 10'hda == io_BankIO_DataAddr ? buffer_218 : _GEN_1241; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1243 = 10'hdb == io_BankIO_DataAddr ? buffer_219 : _GEN_1242; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1244 = 10'hdc == io_BankIO_DataAddr ? buffer_220 : _GEN_1243; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1245 = 10'hdd == io_BankIO_DataAddr ? buffer_221 : _GEN_1244; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1246 = 10'hde == io_BankIO_DataAddr ? buffer_222 : _GEN_1245; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1247 = 10'hdf == io_BankIO_DataAddr ? buffer_223 : _GEN_1246; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1248 = 10'he0 == io_BankIO_DataAddr ? buffer_224 : _GEN_1247; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1249 = 10'he1 == io_BankIO_DataAddr ? buffer_225 : _GEN_1248; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1250 = 10'he2 == io_BankIO_DataAddr ? buffer_226 : _GEN_1249; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1251 = 10'he3 == io_BankIO_DataAddr ? buffer_227 : _GEN_1250; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1252 = 10'he4 == io_BankIO_DataAddr ? buffer_228 : _GEN_1251; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1253 = 10'he5 == io_BankIO_DataAddr ? buffer_229 : _GEN_1252; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1254 = 10'he6 == io_BankIO_DataAddr ? buffer_230 : _GEN_1253; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1255 = 10'he7 == io_BankIO_DataAddr ? buffer_231 : _GEN_1254; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1256 = 10'he8 == io_BankIO_DataAddr ? buffer_232 : _GEN_1255; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1257 = 10'he9 == io_BankIO_DataAddr ? buffer_233 : _GEN_1256; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1258 = 10'hea == io_BankIO_DataAddr ? buffer_234 : _GEN_1257; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1259 = 10'heb == io_BankIO_DataAddr ? buffer_235 : _GEN_1258; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1260 = 10'hec == io_BankIO_DataAddr ? buffer_236 : _GEN_1259; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1261 = 10'hed == io_BankIO_DataAddr ? buffer_237 : _GEN_1260; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1262 = 10'hee == io_BankIO_DataAddr ? buffer_238 : _GEN_1261; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1263 = 10'hef == io_BankIO_DataAddr ? buffer_239 : _GEN_1262; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1264 = 10'hf0 == io_BankIO_DataAddr ? buffer_240 : _GEN_1263; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1265 = 10'hf1 == io_BankIO_DataAddr ? buffer_241 : _GEN_1264; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1266 = 10'hf2 == io_BankIO_DataAddr ? buffer_242 : _GEN_1265; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1267 = 10'hf3 == io_BankIO_DataAddr ? buffer_243 : _GEN_1266; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1268 = 10'hf4 == io_BankIO_DataAddr ? buffer_244 : _GEN_1267; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1269 = 10'hf5 == io_BankIO_DataAddr ? buffer_245 : _GEN_1268; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1270 = 10'hf6 == io_BankIO_DataAddr ? buffer_246 : _GEN_1269; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1271 = 10'hf7 == io_BankIO_DataAddr ? buffer_247 : _GEN_1270; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1272 = 10'hf8 == io_BankIO_DataAddr ? buffer_248 : _GEN_1271; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1273 = 10'hf9 == io_BankIO_DataAddr ? buffer_249 : _GEN_1272; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1274 = 10'hfa == io_BankIO_DataAddr ? buffer_250 : _GEN_1273; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1275 = 10'hfb == io_BankIO_DataAddr ? buffer_251 : _GEN_1274; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1276 = 10'hfc == io_BankIO_DataAddr ? buffer_252 : _GEN_1275; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1277 = 10'hfd == io_BankIO_DataAddr ? buffer_253 : _GEN_1276; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1278 = 10'hfe == io_BankIO_DataAddr ? buffer_254 : _GEN_1277; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1279 = 10'hff == io_BankIO_DataAddr ? buffer_255 : _GEN_1278; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1280 = 10'h100 == io_BankIO_DataAddr ? buffer_256 : _GEN_1279; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1281 = 10'h101 == io_BankIO_DataAddr ? buffer_257 : _GEN_1280; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1282 = 10'h102 == io_BankIO_DataAddr ? buffer_258 : _GEN_1281; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1283 = 10'h103 == io_BankIO_DataAddr ? buffer_259 : _GEN_1282; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1284 = 10'h104 == io_BankIO_DataAddr ? buffer_260 : _GEN_1283; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1285 = 10'h105 == io_BankIO_DataAddr ? buffer_261 : _GEN_1284; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1286 = 10'h106 == io_BankIO_DataAddr ? buffer_262 : _GEN_1285; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1287 = 10'h107 == io_BankIO_DataAddr ? buffer_263 : _GEN_1286; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1288 = 10'h108 == io_BankIO_DataAddr ? buffer_264 : _GEN_1287; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1289 = 10'h109 == io_BankIO_DataAddr ? buffer_265 : _GEN_1288; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1290 = 10'h10a == io_BankIO_DataAddr ? buffer_266 : _GEN_1289; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1291 = 10'h10b == io_BankIO_DataAddr ? buffer_267 : _GEN_1290; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1292 = 10'h10c == io_BankIO_DataAddr ? buffer_268 : _GEN_1291; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1293 = 10'h10d == io_BankIO_DataAddr ? buffer_269 : _GEN_1292; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1294 = 10'h10e == io_BankIO_DataAddr ? buffer_270 : _GEN_1293; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1295 = 10'h10f == io_BankIO_DataAddr ? buffer_271 : _GEN_1294; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1296 = 10'h110 == io_BankIO_DataAddr ? buffer_272 : _GEN_1295; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1297 = 10'h111 == io_BankIO_DataAddr ? buffer_273 : _GEN_1296; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1298 = 10'h112 == io_BankIO_DataAddr ? buffer_274 : _GEN_1297; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1299 = 10'h113 == io_BankIO_DataAddr ? buffer_275 : _GEN_1298; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1300 = 10'h114 == io_BankIO_DataAddr ? buffer_276 : _GEN_1299; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1301 = 10'h115 == io_BankIO_DataAddr ? buffer_277 : _GEN_1300; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1302 = 10'h116 == io_BankIO_DataAddr ? buffer_278 : _GEN_1301; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1303 = 10'h117 == io_BankIO_DataAddr ? buffer_279 : _GEN_1302; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1304 = 10'h118 == io_BankIO_DataAddr ? buffer_280 : _GEN_1303; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1305 = 10'h119 == io_BankIO_DataAddr ? buffer_281 : _GEN_1304; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1306 = 10'h11a == io_BankIO_DataAddr ? buffer_282 : _GEN_1305; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1307 = 10'h11b == io_BankIO_DataAddr ? buffer_283 : _GEN_1306; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1308 = 10'h11c == io_BankIO_DataAddr ? buffer_284 : _GEN_1307; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1309 = 10'h11d == io_BankIO_DataAddr ? buffer_285 : _GEN_1308; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1310 = 10'h11e == io_BankIO_DataAddr ? buffer_286 : _GEN_1309; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1311 = 10'h11f == io_BankIO_DataAddr ? buffer_287 : _GEN_1310; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1312 = 10'h120 == io_BankIO_DataAddr ? buffer_288 : _GEN_1311; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1313 = 10'h121 == io_BankIO_DataAddr ? buffer_289 : _GEN_1312; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1314 = 10'h122 == io_BankIO_DataAddr ? buffer_290 : _GEN_1313; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1315 = 10'h123 == io_BankIO_DataAddr ? buffer_291 : _GEN_1314; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1316 = 10'h124 == io_BankIO_DataAddr ? buffer_292 : _GEN_1315; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1317 = 10'h125 == io_BankIO_DataAddr ? buffer_293 : _GEN_1316; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1318 = 10'h126 == io_BankIO_DataAddr ? buffer_294 : _GEN_1317; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1319 = 10'h127 == io_BankIO_DataAddr ? buffer_295 : _GEN_1318; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1320 = 10'h128 == io_BankIO_DataAddr ? buffer_296 : _GEN_1319; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1321 = 10'h129 == io_BankIO_DataAddr ? buffer_297 : _GEN_1320; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1322 = 10'h12a == io_BankIO_DataAddr ? buffer_298 : _GEN_1321; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1323 = 10'h12b == io_BankIO_DataAddr ? buffer_299 : _GEN_1322; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1324 = 10'h12c == io_BankIO_DataAddr ? buffer_300 : _GEN_1323; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1325 = 10'h12d == io_BankIO_DataAddr ? buffer_301 : _GEN_1324; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1326 = 10'h12e == io_BankIO_DataAddr ? buffer_302 : _GEN_1325; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1327 = 10'h12f == io_BankIO_DataAddr ? buffer_303 : _GEN_1326; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1328 = 10'h130 == io_BankIO_DataAddr ? buffer_304 : _GEN_1327; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1329 = 10'h131 == io_BankIO_DataAddr ? buffer_305 : _GEN_1328; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1330 = 10'h132 == io_BankIO_DataAddr ? buffer_306 : _GEN_1329; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1331 = 10'h133 == io_BankIO_DataAddr ? buffer_307 : _GEN_1330; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1332 = 10'h134 == io_BankIO_DataAddr ? buffer_308 : _GEN_1331; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1333 = 10'h135 == io_BankIO_DataAddr ? buffer_309 : _GEN_1332; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1334 = 10'h136 == io_BankIO_DataAddr ? buffer_310 : _GEN_1333; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1335 = 10'h137 == io_BankIO_DataAddr ? buffer_311 : _GEN_1334; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1336 = 10'h138 == io_BankIO_DataAddr ? buffer_312 : _GEN_1335; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1337 = 10'h139 == io_BankIO_DataAddr ? buffer_313 : _GEN_1336; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1338 = 10'h13a == io_BankIO_DataAddr ? buffer_314 : _GEN_1337; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1339 = 10'h13b == io_BankIO_DataAddr ? buffer_315 : _GEN_1338; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1340 = 10'h13c == io_BankIO_DataAddr ? buffer_316 : _GEN_1339; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1341 = 10'h13d == io_BankIO_DataAddr ? buffer_317 : _GEN_1340; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1342 = 10'h13e == io_BankIO_DataAddr ? buffer_318 : _GEN_1341; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1343 = 10'h13f == io_BankIO_DataAddr ? buffer_319 : _GEN_1342; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1344 = 10'h140 == io_BankIO_DataAddr ? buffer_320 : _GEN_1343; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1345 = 10'h141 == io_BankIO_DataAddr ? buffer_321 : _GEN_1344; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1346 = 10'h142 == io_BankIO_DataAddr ? buffer_322 : _GEN_1345; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1347 = 10'h143 == io_BankIO_DataAddr ? buffer_323 : _GEN_1346; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1348 = 10'h144 == io_BankIO_DataAddr ? buffer_324 : _GEN_1347; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1349 = 10'h145 == io_BankIO_DataAddr ? buffer_325 : _GEN_1348; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1350 = 10'h146 == io_BankIO_DataAddr ? buffer_326 : _GEN_1349; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1351 = 10'h147 == io_BankIO_DataAddr ? buffer_327 : _GEN_1350; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1352 = 10'h148 == io_BankIO_DataAddr ? buffer_328 : _GEN_1351; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1353 = 10'h149 == io_BankIO_DataAddr ? buffer_329 : _GEN_1352; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1354 = 10'h14a == io_BankIO_DataAddr ? buffer_330 : _GEN_1353; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1355 = 10'h14b == io_BankIO_DataAddr ? buffer_331 : _GEN_1354; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1356 = 10'h14c == io_BankIO_DataAddr ? buffer_332 : _GEN_1355; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1357 = 10'h14d == io_BankIO_DataAddr ? buffer_333 : _GEN_1356; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1358 = 10'h14e == io_BankIO_DataAddr ? buffer_334 : _GEN_1357; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1359 = 10'h14f == io_BankIO_DataAddr ? buffer_335 : _GEN_1358; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1360 = 10'h150 == io_BankIO_DataAddr ? buffer_336 : _GEN_1359; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1361 = 10'h151 == io_BankIO_DataAddr ? buffer_337 : _GEN_1360; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1362 = 10'h152 == io_BankIO_DataAddr ? buffer_338 : _GEN_1361; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1363 = 10'h153 == io_BankIO_DataAddr ? buffer_339 : _GEN_1362; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1364 = 10'h154 == io_BankIO_DataAddr ? buffer_340 : _GEN_1363; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1365 = 10'h155 == io_BankIO_DataAddr ? buffer_341 : _GEN_1364; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1366 = 10'h156 == io_BankIO_DataAddr ? buffer_342 : _GEN_1365; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1367 = 10'h157 == io_BankIO_DataAddr ? buffer_343 : _GEN_1366; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1368 = 10'h158 == io_BankIO_DataAddr ? buffer_344 : _GEN_1367; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1369 = 10'h159 == io_BankIO_DataAddr ? buffer_345 : _GEN_1368; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1370 = 10'h15a == io_BankIO_DataAddr ? buffer_346 : _GEN_1369; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1371 = 10'h15b == io_BankIO_DataAddr ? buffer_347 : _GEN_1370; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1372 = 10'h15c == io_BankIO_DataAddr ? buffer_348 : _GEN_1371; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1373 = 10'h15d == io_BankIO_DataAddr ? buffer_349 : _GEN_1372; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1374 = 10'h15e == io_BankIO_DataAddr ? buffer_350 : _GEN_1373; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1375 = 10'h15f == io_BankIO_DataAddr ? buffer_351 : _GEN_1374; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1376 = 10'h160 == io_BankIO_DataAddr ? buffer_352 : _GEN_1375; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1377 = 10'h161 == io_BankIO_DataAddr ? buffer_353 : _GEN_1376; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1378 = 10'h162 == io_BankIO_DataAddr ? buffer_354 : _GEN_1377; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1379 = 10'h163 == io_BankIO_DataAddr ? buffer_355 : _GEN_1378; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1380 = 10'h164 == io_BankIO_DataAddr ? buffer_356 : _GEN_1379; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1381 = 10'h165 == io_BankIO_DataAddr ? buffer_357 : _GEN_1380; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1382 = 10'h166 == io_BankIO_DataAddr ? buffer_358 : _GEN_1381; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1383 = 10'h167 == io_BankIO_DataAddr ? buffer_359 : _GEN_1382; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1384 = 10'h168 == io_BankIO_DataAddr ? buffer_360 : _GEN_1383; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1385 = 10'h169 == io_BankIO_DataAddr ? buffer_361 : _GEN_1384; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1386 = 10'h16a == io_BankIO_DataAddr ? buffer_362 : _GEN_1385; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1387 = 10'h16b == io_BankIO_DataAddr ? buffer_363 : _GEN_1386; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1388 = 10'h16c == io_BankIO_DataAddr ? buffer_364 : _GEN_1387; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1389 = 10'h16d == io_BankIO_DataAddr ? buffer_365 : _GEN_1388; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1390 = 10'h16e == io_BankIO_DataAddr ? buffer_366 : _GEN_1389; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1391 = 10'h16f == io_BankIO_DataAddr ? buffer_367 : _GEN_1390; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1392 = 10'h170 == io_BankIO_DataAddr ? buffer_368 : _GEN_1391; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1393 = 10'h171 == io_BankIO_DataAddr ? buffer_369 : _GEN_1392; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1394 = 10'h172 == io_BankIO_DataAddr ? buffer_370 : _GEN_1393; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1395 = 10'h173 == io_BankIO_DataAddr ? buffer_371 : _GEN_1394; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1396 = 10'h174 == io_BankIO_DataAddr ? buffer_372 : _GEN_1395; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1397 = 10'h175 == io_BankIO_DataAddr ? buffer_373 : _GEN_1396; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1398 = 10'h176 == io_BankIO_DataAddr ? buffer_374 : _GEN_1397; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1399 = 10'h177 == io_BankIO_DataAddr ? buffer_375 : _GEN_1398; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1400 = 10'h178 == io_BankIO_DataAddr ? buffer_376 : _GEN_1399; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1401 = 10'h179 == io_BankIO_DataAddr ? buffer_377 : _GEN_1400; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1402 = 10'h17a == io_BankIO_DataAddr ? buffer_378 : _GEN_1401; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1403 = 10'h17b == io_BankIO_DataAddr ? buffer_379 : _GEN_1402; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1404 = 10'h17c == io_BankIO_DataAddr ? buffer_380 : _GEN_1403; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1405 = 10'h17d == io_BankIO_DataAddr ? buffer_381 : _GEN_1404; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1406 = 10'h17e == io_BankIO_DataAddr ? buffer_382 : _GEN_1405; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1407 = 10'h17f == io_BankIO_DataAddr ? buffer_383 : _GEN_1406; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1408 = 10'h180 == io_BankIO_DataAddr ? buffer_384 : _GEN_1407; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1409 = 10'h181 == io_BankIO_DataAddr ? buffer_385 : _GEN_1408; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1410 = 10'h182 == io_BankIO_DataAddr ? buffer_386 : _GEN_1409; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1411 = 10'h183 == io_BankIO_DataAddr ? buffer_387 : _GEN_1410; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1412 = 10'h184 == io_BankIO_DataAddr ? buffer_388 : _GEN_1411; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1413 = 10'h185 == io_BankIO_DataAddr ? buffer_389 : _GEN_1412; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1414 = 10'h186 == io_BankIO_DataAddr ? buffer_390 : _GEN_1413; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1415 = 10'h187 == io_BankIO_DataAddr ? buffer_391 : _GEN_1414; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1416 = 10'h188 == io_BankIO_DataAddr ? buffer_392 : _GEN_1415; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1417 = 10'h189 == io_BankIO_DataAddr ? buffer_393 : _GEN_1416; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1418 = 10'h18a == io_BankIO_DataAddr ? buffer_394 : _GEN_1417; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1419 = 10'h18b == io_BankIO_DataAddr ? buffer_395 : _GEN_1418; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1420 = 10'h18c == io_BankIO_DataAddr ? buffer_396 : _GEN_1419; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1421 = 10'h18d == io_BankIO_DataAddr ? buffer_397 : _GEN_1420; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1422 = 10'h18e == io_BankIO_DataAddr ? buffer_398 : _GEN_1421; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1423 = 10'h18f == io_BankIO_DataAddr ? buffer_399 : _GEN_1422; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1424 = 10'h190 == io_BankIO_DataAddr ? buffer_400 : _GEN_1423; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1425 = 10'h191 == io_BankIO_DataAddr ? buffer_401 : _GEN_1424; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1426 = 10'h192 == io_BankIO_DataAddr ? buffer_402 : _GEN_1425; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1427 = 10'h193 == io_BankIO_DataAddr ? buffer_403 : _GEN_1426; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1428 = 10'h194 == io_BankIO_DataAddr ? buffer_404 : _GEN_1427; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1429 = 10'h195 == io_BankIO_DataAddr ? buffer_405 : _GEN_1428; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1430 = 10'h196 == io_BankIO_DataAddr ? buffer_406 : _GEN_1429; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1431 = 10'h197 == io_BankIO_DataAddr ? buffer_407 : _GEN_1430; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1432 = 10'h198 == io_BankIO_DataAddr ? buffer_408 : _GEN_1431; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1433 = 10'h199 == io_BankIO_DataAddr ? buffer_409 : _GEN_1432; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1434 = 10'h19a == io_BankIO_DataAddr ? buffer_410 : _GEN_1433; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1435 = 10'h19b == io_BankIO_DataAddr ? buffer_411 : _GEN_1434; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1436 = 10'h19c == io_BankIO_DataAddr ? buffer_412 : _GEN_1435; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1437 = 10'h19d == io_BankIO_DataAddr ? buffer_413 : _GEN_1436; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1438 = 10'h19e == io_BankIO_DataAddr ? buffer_414 : _GEN_1437; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1439 = 10'h19f == io_BankIO_DataAddr ? buffer_415 : _GEN_1438; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1440 = 10'h1a0 == io_BankIO_DataAddr ? buffer_416 : _GEN_1439; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1441 = 10'h1a1 == io_BankIO_DataAddr ? buffer_417 : _GEN_1440; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1442 = 10'h1a2 == io_BankIO_DataAddr ? buffer_418 : _GEN_1441; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1443 = 10'h1a3 == io_BankIO_DataAddr ? buffer_419 : _GEN_1442; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1444 = 10'h1a4 == io_BankIO_DataAddr ? buffer_420 : _GEN_1443; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1445 = 10'h1a5 == io_BankIO_DataAddr ? buffer_421 : _GEN_1444; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1446 = 10'h1a6 == io_BankIO_DataAddr ? buffer_422 : _GEN_1445; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1447 = 10'h1a7 == io_BankIO_DataAddr ? buffer_423 : _GEN_1446; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1448 = 10'h1a8 == io_BankIO_DataAddr ? buffer_424 : _GEN_1447; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1449 = 10'h1a9 == io_BankIO_DataAddr ? buffer_425 : _GEN_1448; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1450 = 10'h1aa == io_BankIO_DataAddr ? buffer_426 : _GEN_1449; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1451 = 10'h1ab == io_BankIO_DataAddr ? buffer_427 : _GEN_1450; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1452 = 10'h1ac == io_BankIO_DataAddr ? buffer_428 : _GEN_1451; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1453 = 10'h1ad == io_BankIO_DataAddr ? buffer_429 : _GEN_1452; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1454 = 10'h1ae == io_BankIO_DataAddr ? buffer_430 : _GEN_1453; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1455 = 10'h1af == io_BankIO_DataAddr ? buffer_431 : _GEN_1454; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1456 = 10'h1b0 == io_BankIO_DataAddr ? buffer_432 : _GEN_1455; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1457 = 10'h1b1 == io_BankIO_DataAddr ? buffer_433 : _GEN_1456; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1458 = 10'h1b2 == io_BankIO_DataAddr ? buffer_434 : _GEN_1457; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1459 = 10'h1b3 == io_BankIO_DataAddr ? buffer_435 : _GEN_1458; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1460 = 10'h1b4 == io_BankIO_DataAddr ? buffer_436 : _GEN_1459; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1461 = 10'h1b5 == io_BankIO_DataAddr ? buffer_437 : _GEN_1460; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1462 = 10'h1b6 == io_BankIO_DataAddr ? buffer_438 : _GEN_1461; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1463 = 10'h1b7 == io_BankIO_DataAddr ? buffer_439 : _GEN_1462; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1464 = 10'h1b8 == io_BankIO_DataAddr ? buffer_440 : _GEN_1463; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1465 = 10'h1b9 == io_BankIO_DataAddr ? buffer_441 : _GEN_1464; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1466 = 10'h1ba == io_BankIO_DataAddr ? buffer_442 : _GEN_1465; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1467 = 10'h1bb == io_BankIO_DataAddr ? buffer_443 : _GEN_1466; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1468 = 10'h1bc == io_BankIO_DataAddr ? buffer_444 : _GEN_1467; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1469 = 10'h1bd == io_BankIO_DataAddr ? buffer_445 : _GEN_1468; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1470 = 10'h1be == io_BankIO_DataAddr ? buffer_446 : _GEN_1469; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1471 = 10'h1bf == io_BankIO_DataAddr ? buffer_447 : _GEN_1470; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1472 = 10'h1c0 == io_BankIO_DataAddr ? buffer_448 : _GEN_1471; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1473 = 10'h1c1 == io_BankIO_DataAddr ? buffer_449 : _GEN_1472; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1474 = 10'h1c2 == io_BankIO_DataAddr ? buffer_450 : _GEN_1473; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1475 = 10'h1c3 == io_BankIO_DataAddr ? buffer_451 : _GEN_1474; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1476 = 10'h1c4 == io_BankIO_DataAddr ? buffer_452 : _GEN_1475; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1477 = 10'h1c5 == io_BankIO_DataAddr ? buffer_453 : _GEN_1476; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1478 = 10'h1c6 == io_BankIO_DataAddr ? buffer_454 : _GEN_1477; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1479 = 10'h1c7 == io_BankIO_DataAddr ? buffer_455 : _GEN_1478; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1480 = 10'h1c8 == io_BankIO_DataAddr ? buffer_456 : _GEN_1479; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1481 = 10'h1c9 == io_BankIO_DataAddr ? buffer_457 : _GEN_1480; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1482 = 10'h1ca == io_BankIO_DataAddr ? buffer_458 : _GEN_1481; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1483 = 10'h1cb == io_BankIO_DataAddr ? buffer_459 : _GEN_1482; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1484 = 10'h1cc == io_BankIO_DataAddr ? buffer_460 : _GEN_1483; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1485 = 10'h1cd == io_BankIO_DataAddr ? buffer_461 : _GEN_1484; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1486 = 10'h1ce == io_BankIO_DataAddr ? buffer_462 : _GEN_1485; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1487 = 10'h1cf == io_BankIO_DataAddr ? buffer_463 : _GEN_1486; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1488 = 10'h1d0 == io_BankIO_DataAddr ? buffer_464 : _GEN_1487; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1489 = 10'h1d1 == io_BankIO_DataAddr ? buffer_465 : _GEN_1488; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1490 = 10'h1d2 == io_BankIO_DataAddr ? buffer_466 : _GEN_1489; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1491 = 10'h1d3 == io_BankIO_DataAddr ? buffer_467 : _GEN_1490; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1492 = 10'h1d4 == io_BankIO_DataAddr ? buffer_468 : _GEN_1491; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1493 = 10'h1d5 == io_BankIO_DataAddr ? buffer_469 : _GEN_1492; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1494 = 10'h1d6 == io_BankIO_DataAddr ? buffer_470 : _GEN_1493; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1495 = 10'h1d7 == io_BankIO_DataAddr ? buffer_471 : _GEN_1494; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1496 = 10'h1d8 == io_BankIO_DataAddr ? buffer_472 : _GEN_1495; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1497 = 10'h1d9 == io_BankIO_DataAddr ? buffer_473 : _GEN_1496; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1498 = 10'h1da == io_BankIO_DataAddr ? buffer_474 : _GEN_1497; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1499 = 10'h1db == io_BankIO_DataAddr ? buffer_475 : _GEN_1498; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1500 = 10'h1dc == io_BankIO_DataAddr ? buffer_476 : _GEN_1499; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1501 = 10'h1dd == io_BankIO_DataAddr ? buffer_477 : _GEN_1500; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1502 = 10'h1de == io_BankIO_DataAddr ? buffer_478 : _GEN_1501; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1503 = 10'h1df == io_BankIO_DataAddr ? buffer_479 : _GEN_1502; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1504 = 10'h1e0 == io_BankIO_DataAddr ? buffer_480 : _GEN_1503; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1505 = 10'h1e1 == io_BankIO_DataAddr ? buffer_481 : _GEN_1504; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1506 = 10'h1e2 == io_BankIO_DataAddr ? buffer_482 : _GEN_1505; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1507 = 10'h1e3 == io_BankIO_DataAddr ? buffer_483 : _GEN_1506; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1508 = 10'h1e4 == io_BankIO_DataAddr ? buffer_484 : _GEN_1507; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1509 = 10'h1e5 == io_BankIO_DataAddr ? buffer_485 : _GEN_1508; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1510 = 10'h1e6 == io_BankIO_DataAddr ? buffer_486 : _GEN_1509; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1511 = 10'h1e7 == io_BankIO_DataAddr ? buffer_487 : _GEN_1510; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1512 = 10'h1e8 == io_BankIO_DataAddr ? buffer_488 : _GEN_1511; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1513 = 10'h1e9 == io_BankIO_DataAddr ? buffer_489 : _GEN_1512; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1514 = 10'h1ea == io_BankIO_DataAddr ? buffer_490 : _GEN_1513; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1515 = 10'h1eb == io_BankIO_DataAddr ? buffer_491 : _GEN_1514; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1516 = 10'h1ec == io_BankIO_DataAddr ? buffer_492 : _GEN_1515; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1517 = 10'h1ed == io_BankIO_DataAddr ? buffer_493 : _GEN_1516; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1518 = 10'h1ee == io_BankIO_DataAddr ? buffer_494 : _GEN_1517; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1519 = 10'h1ef == io_BankIO_DataAddr ? buffer_495 : _GEN_1518; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1520 = 10'h1f0 == io_BankIO_DataAddr ? buffer_496 : _GEN_1519; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1521 = 10'h1f1 == io_BankIO_DataAddr ? buffer_497 : _GEN_1520; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1522 = 10'h1f2 == io_BankIO_DataAddr ? buffer_498 : _GEN_1521; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1523 = 10'h1f3 == io_BankIO_DataAddr ? buffer_499 : _GEN_1522; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1524 = 10'h1f4 == io_BankIO_DataAddr ? buffer_500 : _GEN_1523; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1525 = 10'h1f5 == io_BankIO_DataAddr ? buffer_501 : _GEN_1524; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1526 = 10'h1f6 == io_BankIO_DataAddr ? buffer_502 : _GEN_1525; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1527 = 10'h1f7 == io_BankIO_DataAddr ? buffer_503 : _GEN_1526; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1528 = 10'h1f8 == io_BankIO_DataAddr ? buffer_504 : _GEN_1527; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1529 = 10'h1f9 == io_BankIO_DataAddr ? buffer_505 : _GEN_1528; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1530 = 10'h1fa == io_BankIO_DataAddr ? buffer_506 : _GEN_1529; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1531 = 10'h1fb == io_BankIO_DataAddr ? buffer_507 : _GEN_1530; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1532 = 10'h1fc == io_BankIO_DataAddr ? buffer_508 : _GEN_1531; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1533 = 10'h1fd == io_BankIO_DataAddr ? buffer_509 : _GEN_1532; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1534 = 10'h1fe == io_BankIO_DataAddr ? buffer_510 : _GEN_1533; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1535 = 10'h1ff == io_BankIO_DataAddr ? buffer_511 : _GEN_1534; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1536 = 10'h200 == io_BankIO_DataAddr ? buffer_512 : _GEN_1535; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1537 = 10'h201 == io_BankIO_DataAddr ? buffer_513 : _GEN_1536; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1538 = 10'h202 == io_BankIO_DataAddr ? buffer_514 : _GEN_1537; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1539 = 10'h203 == io_BankIO_DataAddr ? buffer_515 : _GEN_1538; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1540 = 10'h204 == io_BankIO_DataAddr ? buffer_516 : _GEN_1539; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1541 = 10'h205 == io_BankIO_DataAddr ? buffer_517 : _GEN_1540; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1542 = 10'h206 == io_BankIO_DataAddr ? buffer_518 : _GEN_1541; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1543 = 10'h207 == io_BankIO_DataAddr ? buffer_519 : _GEN_1542; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1544 = 10'h208 == io_BankIO_DataAddr ? buffer_520 : _GEN_1543; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1545 = 10'h209 == io_BankIO_DataAddr ? buffer_521 : _GEN_1544; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1546 = 10'h20a == io_BankIO_DataAddr ? buffer_522 : _GEN_1545; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1547 = 10'h20b == io_BankIO_DataAddr ? buffer_523 : _GEN_1546; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1548 = 10'h20c == io_BankIO_DataAddr ? buffer_524 : _GEN_1547; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1549 = 10'h20d == io_BankIO_DataAddr ? buffer_525 : _GEN_1548; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1550 = 10'h20e == io_BankIO_DataAddr ? buffer_526 : _GEN_1549; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1551 = 10'h20f == io_BankIO_DataAddr ? buffer_527 : _GEN_1550; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1552 = 10'h210 == io_BankIO_DataAddr ? buffer_528 : _GEN_1551; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1553 = 10'h211 == io_BankIO_DataAddr ? buffer_529 : _GEN_1552; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1554 = 10'h212 == io_BankIO_DataAddr ? buffer_530 : _GEN_1553; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1555 = 10'h213 == io_BankIO_DataAddr ? buffer_531 : _GEN_1554; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1556 = 10'h214 == io_BankIO_DataAddr ? buffer_532 : _GEN_1555; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1557 = 10'h215 == io_BankIO_DataAddr ? buffer_533 : _GEN_1556; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1558 = 10'h216 == io_BankIO_DataAddr ? buffer_534 : _GEN_1557; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1559 = 10'h217 == io_BankIO_DataAddr ? buffer_535 : _GEN_1558; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1560 = 10'h218 == io_BankIO_DataAddr ? buffer_536 : _GEN_1559; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1561 = 10'h219 == io_BankIO_DataAddr ? buffer_537 : _GEN_1560; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1562 = 10'h21a == io_BankIO_DataAddr ? buffer_538 : _GEN_1561; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1563 = 10'h21b == io_BankIO_DataAddr ? buffer_539 : _GEN_1562; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1564 = 10'h21c == io_BankIO_DataAddr ? buffer_540 : _GEN_1563; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1565 = 10'h21d == io_BankIO_DataAddr ? buffer_541 : _GEN_1564; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1566 = 10'h21e == io_BankIO_DataAddr ? buffer_542 : _GEN_1565; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1567 = 10'h21f == io_BankIO_DataAddr ? buffer_543 : _GEN_1566; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1568 = 10'h220 == io_BankIO_DataAddr ? buffer_544 : _GEN_1567; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1569 = 10'h221 == io_BankIO_DataAddr ? buffer_545 : _GEN_1568; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1570 = 10'h222 == io_BankIO_DataAddr ? buffer_546 : _GEN_1569; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1571 = 10'h223 == io_BankIO_DataAddr ? buffer_547 : _GEN_1570; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1572 = 10'h224 == io_BankIO_DataAddr ? buffer_548 : _GEN_1571; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1573 = 10'h225 == io_BankIO_DataAddr ? buffer_549 : _GEN_1572; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1574 = 10'h226 == io_BankIO_DataAddr ? buffer_550 : _GEN_1573; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1575 = 10'h227 == io_BankIO_DataAddr ? buffer_551 : _GEN_1574; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1576 = 10'h228 == io_BankIO_DataAddr ? buffer_552 : _GEN_1575; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1577 = 10'h229 == io_BankIO_DataAddr ? buffer_553 : _GEN_1576; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1578 = 10'h22a == io_BankIO_DataAddr ? buffer_554 : _GEN_1577; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1579 = 10'h22b == io_BankIO_DataAddr ? buffer_555 : _GEN_1578; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1580 = 10'h22c == io_BankIO_DataAddr ? buffer_556 : _GEN_1579; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1581 = 10'h22d == io_BankIO_DataAddr ? buffer_557 : _GEN_1580; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1582 = 10'h22e == io_BankIO_DataAddr ? buffer_558 : _GEN_1581; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1583 = 10'h22f == io_BankIO_DataAddr ? buffer_559 : _GEN_1582; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1584 = 10'h230 == io_BankIO_DataAddr ? buffer_560 : _GEN_1583; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1585 = 10'h231 == io_BankIO_DataAddr ? buffer_561 : _GEN_1584; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1586 = 10'h232 == io_BankIO_DataAddr ? buffer_562 : _GEN_1585; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1587 = 10'h233 == io_BankIO_DataAddr ? buffer_563 : _GEN_1586; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1588 = 10'h234 == io_BankIO_DataAddr ? buffer_564 : _GEN_1587; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1589 = 10'h235 == io_BankIO_DataAddr ? buffer_565 : _GEN_1588; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1590 = 10'h236 == io_BankIO_DataAddr ? buffer_566 : _GEN_1589; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1591 = 10'h237 == io_BankIO_DataAddr ? buffer_567 : _GEN_1590; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1592 = 10'h238 == io_BankIO_DataAddr ? buffer_568 : _GEN_1591; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1593 = 10'h239 == io_BankIO_DataAddr ? buffer_569 : _GEN_1592; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1594 = 10'h23a == io_BankIO_DataAddr ? buffer_570 : _GEN_1593; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1595 = 10'h23b == io_BankIO_DataAddr ? buffer_571 : _GEN_1594; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1596 = 10'h23c == io_BankIO_DataAddr ? buffer_572 : _GEN_1595; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1597 = 10'h23d == io_BankIO_DataAddr ? buffer_573 : _GEN_1596; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1598 = 10'h23e == io_BankIO_DataAddr ? buffer_574 : _GEN_1597; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1599 = 10'h23f == io_BankIO_DataAddr ? buffer_575 : _GEN_1598; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1600 = 10'h240 == io_BankIO_DataAddr ? buffer_576 : _GEN_1599; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1601 = 10'h241 == io_BankIO_DataAddr ? buffer_577 : _GEN_1600; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1602 = 10'h242 == io_BankIO_DataAddr ? buffer_578 : _GEN_1601; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1603 = 10'h243 == io_BankIO_DataAddr ? buffer_579 : _GEN_1602; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1604 = 10'h244 == io_BankIO_DataAddr ? buffer_580 : _GEN_1603; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1605 = 10'h245 == io_BankIO_DataAddr ? buffer_581 : _GEN_1604; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1606 = 10'h246 == io_BankIO_DataAddr ? buffer_582 : _GEN_1605; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1607 = 10'h247 == io_BankIO_DataAddr ? buffer_583 : _GEN_1606; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1608 = 10'h248 == io_BankIO_DataAddr ? buffer_584 : _GEN_1607; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1609 = 10'h249 == io_BankIO_DataAddr ? buffer_585 : _GEN_1608; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1610 = 10'h24a == io_BankIO_DataAddr ? buffer_586 : _GEN_1609; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1611 = 10'h24b == io_BankIO_DataAddr ? buffer_587 : _GEN_1610; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1612 = 10'h24c == io_BankIO_DataAddr ? buffer_588 : _GEN_1611; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1613 = 10'h24d == io_BankIO_DataAddr ? buffer_589 : _GEN_1612; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1614 = 10'h24e == io_BankIO_DataAddr ? buffer_590 : _GEN_1613; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1615 = 10'h24f == io_BankIO_DataAddr ? buffer_591 : _GEN_1614; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1616 = 10'h250 == io_BankIO_DataAddr ? buffer_592 : _GEN_1615; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1617 = 10'h251 == io_BankIO_DataAddr ? buffer_593 : _GEN_1616; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1618 = 10'h252 == io_BankIO_DataAddr ? buffer_594 : _GEN_1617; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1619 = 10'h253 == io_BankIO_DataAddr ? buffer_595 : _GEN_1618; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1620 = 10'h254 == io_BankIO_DataAddr ? buffer_596 : _GEN_1619; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1621 = 10'h255 == io_BankIO_DataAddr ? buffer_597 : _GEN_1620; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1622 = 10'h256 == io_BankIO_DataAddr ? buffer_598 : _GEN_1621; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1623 = 10'h257 == io_BankIO_DataAddr ? buffer_599 : _GEN_1622; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1624 = 10'h258 == io_BankIO_DataAddr ? buffer_600 : _GEN_1623; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1625 = 10'h259 == io_BankIO_DataAddr ? buffer_601 : _GEN_1624; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1626 = 10'h25a == io_BankIO_DataAddr ? buffer_602 : _GEN_1625; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1627 = 10'h25b == io_BankIO_DataAddr ? buffer_603 : _GEN_1626; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1628 = 10'h25c == io_BankIO_DataAddr ? buffer_604 : _GEN_1627; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1629 = 10'h25d == io_BankIO_DataAddr ? buffer_605 : _GEN_1628; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1630 = 10'h25e == io_BankIO_DataAddr ? buffer_606 : _GEN_1629; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1631 = 10'h25f == io_BankIO_DataAddr ? buffer_607 : _GEN_1630; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1632 = 10'h260 == io_BankIO_DataAddr ? buffer_608 : _GEN_1631; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1633 = 10'h261 == io_BankIO_DataAddr ? buffer_609 : _GEN_1632; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1634 = 10'h262 == io_BankIO_DataAddr ? buffer_610 : _GEN_1633; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1635 = 10'h263 == io_BankIO_DataAddr ? buffer_611 : _GEN_1634; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1636 = 10'h264 == io_BankIO_DataAddr ? buffer_612 : _GEN_1635; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1637 = 10'h265 == io_BankIO_DataAddr ? buffer_613 : _GEN_1636; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1638 = 10'h266 == io_BankIO_DataAddr ? buffer_614 : _GEN_1637; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1639 = 10'h267 == io_BankIO_DataAddr ? buffer_615 : _GEN_1638; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1640 = 10'h268 == io_BankIO_DataAddr ? buffer_616 : _GEN_1639; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1641 = 10'h269 == io_BankIO_DataAddr ? buffer_617 : _GEN_1640; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1642 = 10'h26a == io_BankIO_DataAddr ? buffer_618 : _GEN_1641; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1643 = 10'h26b == io_BankIO_DataAddr ? buffer_619 : _GEN_1642; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1644 = 10'h26c == io_BankIO_DataAddr ? buffer_620 : _GEN_1643; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1645 = 10'h26d == io_BankIO_DataAddr ? buffer_621 : _GEN_1644; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1646 = 10'h26e == io_BankIO_DataAddr ? buffer_622 : _GEN_1645; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1647 = 10'h26f == io_BankIO_DataAddr ? buffer_623 : _GEN_1646; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1648 = 10'h270 == io_BankIO_DataAddr ? buffer_624 : _GEN_1647; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1649 = 10'h271 == io_BankIO_DataAddr ? buffer_625 : _GEN_1648; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1650 = 10'h272 == io_BankIO_DataAddr ? buffer_626 : _GEN_1649; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1651 = 10'h273 == io_BankIO_DataAddr ? buffer_627 : _GEN_1650; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1652 = 10'h274 == io_BankIO_DataAddr ? buffer_628 : _GEN_1651; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1653 = 10'h275 == io_BankIO_DataAddr ? buffer_629 : _GEN_1652; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1654 = 10'h276 == io_BankIO_DataAddr ? buffer_630 : _GEN_1653; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1655 = 10'h277 == io_BankIO_DataAddr ? buffer_631 : _GEN_1654; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1656 = 10'h278 == io_BankIO_DataAddr ? buffer_632 : _GEN_1655; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1657 = 10'h279 == io_BankIO_DataAddr ? buffer_633 : _GEN_1656; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1658 = 10'h27a == io_BankIO_DataAddr ? buffer_634 : _GEN_1657; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1659 = 10'h27b == io_BankIO_DataAddr ? buffer_635 : _GEN_1658; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1660 = 10'h27c == io_BankIO_DataAddr ? buffer_636 : _GEN_1659; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1661 = 10'h27d == io_BankIO_DataAddr ? buffer_637 : _GEN_1660; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1662 = 10'h27e == io_BankIO_DataAddr ? buffer_638 : _GEN_1661; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1663 = 10'h27f == io_BankIO_DataAddr ? buffer_639 : _GEN_1662; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1664 = 10'h280 == io_BankIO_DataAddr ? buffer_640 : _GEN_1663; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1665 = 10'h281 == io_BankIO_DataAddr ? buffer_641 : _GEN_1664; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1666 = 10'h282 == io_BankIO_DataAddr ? buffer_642 : _GEN_1665; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1667 = 10'h283 == io_BankIO_DataAddr ? buffer_643 : _GEN_1666; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1668 = 10'h284 == io_BankIO_DataAddr ? buffer_644 : _GEN_1667; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1669 = 10'h285 == io_BankIO_DataAddr ? buffer_645 : _GEN_1668; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1670 = 10'h286 == io_BankIO_DataAddr ? buffer_646 : _GEN_1669; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1671 = 10'h287 == io_BankIO_DataAddr ? buffer_647 : _GEN_1670; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1672 = 10'h288 == io_BankIO_DataAddr ? buffer_648 : _GEN_1671; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1673 = 10'h289 == io_BankIO_DataAddr ? buffer_649 : _GEN_1672; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1674 = 10'h28a == io_BankIO_DataAddr ? buffer_650 : _GEN_1673; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1675 = 10'h28b == io_BankIO_DataAddr ? buffer_651 : _GEN_1674; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1676 = 10'h28c == io_BankIO_DataAddr ? buffer_652 : _GEN_1675; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1677 = 10'h28d == io_BankIO_DataAddr ? buffer_653 : _GEN_1676; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1678 = 10'h28e == io_BankIO_DataAddr ? buffer_654 : _GEN_1677; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1679 = 10'h28f == io_BankIO_DataAddr ? buffer_655 : _GEN_1678; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1680 = 10'h290 == io_BankIO_DataAddr ? buffer_656 : _GEN_1679; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1681 = 10'h291 == io_BankIO_DataAddr ? buffer_657 : _GEN_1680; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1682 = 10'h292 == io_BankIO_DataAddr ? buffer_658 : _GEN_1681; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1683 = 10'h293 == io_BankIO_DataAddr ? buffer_659 : _GEN_1682; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1684 = 10'h294 == io_BankIO_DataAddr ? buffer_660 : _GEN_1683; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1685 = 10'h295 == io_BankIO_DataAddr ? buffer_661 : _GEN_1684; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1686 = 10'h296 == io_BankIO_DataAddr ? buffer_662 : _GEN_1685; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1687 = 10'h297 == io_BankIO_DataAddr ? buffer_663 : _GEN_1686; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1688 = 10'h298 == io_BankIO_DataAddr ? buffer_664 : _GEN_1687; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1689 = 10'h299 == io_BankIO_DataAddr ? buffer_665 : _GEN_1688; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1690 = 10'h29a == io_BankIO_DataAddr ? buffer_666 : _GEN_1689; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1691 = 10'h29b == io_BankIO_DataAddr ? buffer_667 : _GEN_1690; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1692 = 10'h29c == io_BankIO_DataAddr ? buffer_668 : _GEN_1691; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1693 = 10'h29d == io_BankIO_DataAddr ? buffer_669 : _GEN_1692; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1694 = 10'h29e == io_BankIO_DataAddr ? buffer_670 : _GEN_1693; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1695 = 10'h29f == io_BankIO_DataAddr ? buffer_671 : _GEN_1694; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1696 = 10'h2a0 == io_BankIO_DataAddr ? buffer_672 : _GEN_1695; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1697 = 10'h2a1 == io_BankIO_DataAddr ? buffer_673 : _GEN_1696; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1698 = 10'h2a2 == io_BankIO_DataAddr ? buffer_674 : _GEN_1697; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1699 = 10'h2a3 == io_BankIO_DataAddr ? buffer_675 : _GEN_1698; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1700 = 10'h2a4 == io_BankIO_DataAddr ? buffer_676 : _GEN_1699; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1701 = 10'h2a5 == io_BankIO_DataAddr ? buffer_677 : _GEN_1700; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1702 = 10'h2a6 == io_BankIO_DataAddr ? buffer_678 : _GEN_1701; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1703 = 10'h2a7 == io_BankIO_DataAddr ? buffer_679 : _GEN_1702; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1704 = 10'h2a8 == io_BankIO_DataAddr ? buffer_680 : _GEN_1703; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1705 = 10'h2a9 == io_BankIO_DataAddr ? buffer_681 : _GEN_1704; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1706 = 10'h2aa == io_BankIO_DataAddr ? buffer_682 : _GEN_1705; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1707 = 10'h2ab == io_BankIO_DataAddr ? buffer_683 : _GEN_1706; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1708 = 10'h2ac == io_BankIO_DataAddr ? buffer_684 : _GEN_1707; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1709 = 10'h2ad == io_BankIO_DataAddr ? buffer_685 : _GEN_1708; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1710 = 10'h2ae == io_BankIO_DataAddr ? buffer_686 : _GEN_1709; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1711 = 10'h2af == io_BankIO_DataAddr ? buffer_687 : _GEN_1710; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1712 = 10'h2b0 == io_BankIO_DataAddr ? buffer_688 : _GEN_1711; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1713 = 10'h2b1 == io_BankIO_DataAddr ? buffer_689 : _GEN_1712; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1714 = 10'h2b2 == io_BankIO_DataAddr ? buffer_690 : _GEN_1713; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1715 = 10'h2b3 == io_BankIO_DataAddr ? buffer_691 : _GEN_1714; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1716 = 10'h2b4 == io_BankIO_DataAddr ? buffer_692 : _GEN_1715; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1717 = 10'h2b5 == io_BankIO_DataAddr ? buffer_693 : _GEN_1716; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1718 = 10'h2b6 == io_BankIO_DataAddr ? buffer_694 : _GEN_1717; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1719 = 10'h2b7 == io_BankIO_DataAddr ? buffer_695 : _GEN_1718; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1720 = 10'h2b8 == io_BankIO_DataAddr ? buffer_696 : _GEN_1719; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1721 = 10'h2b9 == io_BankIO_DataAddr ? buffer_697 : _GEN_1720; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1722 = 10'h2ba == io_BankIO_DataAddr ? buffer_698 : _GEN_1721; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1723 = 10'h2bb == io_BankIO_DataAddr ? buffer_699 : _GEN_1722; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1724 = 10'h2bc == io_BankIO_DataAddr ? buffer_700 : _GEN_1723; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1725 = 10'h2bd == io_BankIO_DataAddr ? buffer_701 : _GEN_1724; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1726 = 10'h2be == io_BankIO_DataAddr ? buffer_702 : _GEN_1725; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1727 = 10'h2bf == io_BankIO_DataAddr ? buffer_703 : _GEN_1726; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1728 = 10'h2c0 == io_BankIO_DataAddr ? buffer_704 : _GEN_1727; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1729 = 10'h2c1 == io_BankIO_DataAddr ? buffer_705 : _GEN_1728; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1730 = 10'h2c2 == io_BankIO_DataAddr ? buffer_706 : _GEN_1729; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1731 = 10'h2c3 == io_BankIO_DataAddr ? buffer_707 : _GEN_1730; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1732 = 10'h2c4 == io_BankIO_DataAddr ? buffer_708 : _GEN_1731; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1733 = 10'h2c5 == io_BankIO_DataAddr ? buffer_709 : _GEN_1732; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1734 = 10'h2c6 == io_BankIO_DataAddr ? buffer_710 : _GEN_1733; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1735 = 10'h2c7 == io_BankIO_DataAddr ? buffer_711 : _GEN_1734; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1736 = 10'h2c8 == io_BankIO_DataAddr ? buffer_712 : _GEN_1735; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1737 = 10'h2c9 == io_BankIO_DataAddr ? buffer_713 : _GEN_1736; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1738 = 10'h2ca == io_BankIO_DataAddr ? buffer_714 : _GEN_1737; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1739 = 10'h2cb == io_BankIO_DataAddr ? buffer_715 : _GEN_1738; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1740 = 10'h2cc == io_BankIO_DataAddr ? buffer_716 : _GEN_1739; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1741 = 10'h2cd == io_BankIO_DataAddr ? buffer_717 : _GEN_1740; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1742 = 10'h2ce == io_BankIO_DataAddr ? buffer_718 : _GEN_1741; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1743 = 10'h2cf == io_BankIO_DataAddr ? buffer_719 : _GEN_1742; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1744 = 10'h2d0 == io_BankIO_DataAddr ? buffer_720 : _GEN_1743; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1745 = 10'h2d1 == io_BankIO_DataAddr ? buffer_721 : _GEN_1744; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1746 = 10'h2d2 == io_BankIO_DataAddr ? buffer_722 : _GEN_1745; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1747 = 10'h2d3 == io_BankIO_DataAddr ? buffer_723 : _GEN_1746; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1748 = 10'h2d4 == io_BankIO_DataAddr ? buffer_724 : _GEN_1747; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1749 = 10'h2d5 == io_BankIO_DataAddr ? buffer_725 : _GEN_1748; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1750 = 10'h2d6 == io_BankIO_DataAddr ? buffer_726 : _GEN_1749; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1751 = 10'h2d7 == io_BankIO_DataAddr ? buffer_727 : _GEN_1750; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1752 = 10'h2d8 == io_BankIO_DataAddr ? buffer_728 : _GEN_1751; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1753 = 10'h2d9 == io_BankIO_DataAddr ? buffer_729 : _GEN_1752; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1754 = 10'h2da == io_BankIO_DataAddr ? buffer_730 : _GEN_1753; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1755 = 10'h2db == io_BankIO_DataAddr ? buffer_731 : _GEN_1754; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1756 = 10'h2dc == io_BankIO_DataAddr ? buffer_732 : _GEN_1755; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1757 = 10'h2dd == io_BankIO_DataAddr ? buffer_733 : _GEN_1756; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1758 = 10'h2de == io_BankIO_DataAddr ? buffer_734 : _GEN_1757; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1759 = 10'h2df == io_BankIO_DataAddr ? buffer_735 : _GEN_1758; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1760 = 10'h2e0 == io_BankIO_DataAddr ? buffer_736 : _GEN_1759; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1761 = 10'h2e1 == io_BankIO_DataAddr ? buffer_737 : _GEN_1760; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1762 = 10'h2e2 == io_BankIO_DataAddr ? buffer_738 : _GEN_1761; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1763 = 10'h2e3 == io_BankIO_DataAddr ? buffer_739 : _GEN_1762; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1764 = 10'h2e4 == io_BankIO_DataAddr ? buffer_740 : _GEN_1763; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1765 = 10'h2e5 == io_BankIO_DataAddr ? buffer_741 : _GEN_1764; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1766 = 10'h2e6 == io_BankIO_DataAddr ? buffer_742 : _GEN_1765; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1767 = 10'h2e7 == io_BankIO_DataAddr ? buffer_743 : _GEN_1766; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1768 = 10'h2e8 == io_BankIO_DataAddr ? buffer_744 : _GEN_1767; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1769 = 10'h2e9 == io_BankIO_DataAddr ? buffer_745 : _GEN_1768; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1770 = 10'h2ea == io_BankIO_DataAddr ? buffer_746 : _GEN_1769; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1771 = 10'h2eb == io_BankIO_DataAddr ? buffer_747 : _GEN_1770; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1772 = 10'h2ec == io_BankIO_DataAddr ? buffer_748 : _GEN_1771; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1773 = 10'h2ed == io_BankIO_DataAddr ? buffer_749 : _GEN_1772; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1774 = 10'h2ee == io_BankIO_DataAddr ? buffer_750 : _GEN_1773; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1775 = 10'h2ef == io_BankIO_DataAddr ? buffer_751 : _GEN_1774; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1776 = 10'h2f0 == io_BankIO_DataAddr ? buffer_752 : _GEN_1775; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1777 = 10'h2f1 == io_BankIO_DataAddr ? buffer_753 : _GEN_1776; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1778 = 10'h2f2 == io_BankIO_DataAddr ? buffer_754 : _GEN_1777; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1779 = 10'h2f3 == io_BankIO_DataAddr ? buffer_755 : _GEN_1778; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1780 = 10'h2f4 == io_BankIO_DataAddr ? buffer_756 : _GEN_1779; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1781 = 10'h2f5 == io_BankIO_DataAddr ? buffer_757 : _GEN_1780; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1782 = 10'h2f6 == io_BankIO_DataAddr ? buffer_758 : _GEN_1781; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1783 = 10'h2f7 == io_BankIO_DataAddr ? buffer_759 : _GEN_1782; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1784 = 10'h2f8 == io_BankIO_DataAddr ? buffer_760 : _GEN_1783; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1785 = 10'h2f9 == io_BankIO_DataAddr ? buffer_761 : _GEN_1784; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1786 = 10'h2fa == io_BankIO_DataAddr ? buffer_762 : _GEN_1785; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1787 = 10'h2fb == io_BankIO_DataAddr ? buffer_763 : _GEN_1786; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1788 = 10'h2fc == io_BankIO_DataAddr ? buffer_764 : _GEN_1787; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1789 = 10'h2fd == io_BankIO_DataAddr ? buffer_765 : _GEN_1788; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1790 = 10'h2fe == io_BankIO_DataAddr ? buffer_766 : _GEN_1789; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1791 = 10'h2ff == io_BankIO_DataAddr ? buffer_767 : _GEN_1790; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1792 = 10'h300 == io_BankIO_DataAddr ? buffer_768 : _GEN_1791; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1793 = 10'h301 == io_BankIO_DataAddr ? buffer_769 : _GEN_1792; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1794 = 10'h302 == io_BankIO_DataAddr ? buffer_770 : _GEN_1793; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1795 = 10'h303 == io_BankIO_DataAddr ? buffer_771 : _GEN_1794; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1796 = 10'h304 == io_BankIO_DataAddr ? buffer_772 : _GEN_1795; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1797 = 10'h305 == io_BankIO_DataAddr ? buffer_773 : _GEN_1796; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1798 = 10'h306 == io_BankIO_DataAddr ? buffer_774 : _GEN_1797; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1799 = 10'h307 == io_BankIO_DataAddr ? buffer_775 : _GEN_1798; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1800 = 10'h308 == io_BankIO_DataAddr ? buffer_776 : _GEN_1799; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1801 = 10'h309 == io_BankIO_DataAddr ? buffer_777 : _GEN_1800; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1802 = 10'h30a == io_BankIO_DataAddr ? buffer_778 : _GEN_1801; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1803 = 10'h30b == io_BankIO_DataAddr ? buffer_779 : _GEN_1802; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1804 = 10'h30c == io_BankIO_DataAddr ? buffer_780 : _GEN_1803; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1805 = 10'h30d == io_BankIO_DataAddr ? buffer_781 : _GEN_1804; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1806 = 10'h30e == io_BankIO_DataAddr ? buffer_782 : _GEN_1805; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1807 = 10'h30f == io_BankIO_DataAddr ? buffer_783 : _GEN_1806; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1808 = 10'h310 == io_BankIO_DataAddr ? buffer_784 : _GEN_1807; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1809 = 10'h311 == io_BankIO_DataAddr ? buffer_785 : _GEN_1808; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1810 = 10'h312 == io_BankIO_DataAddr ? buffer_786 : _GEN_1809; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1811 = 10'h313 == io_BankIO_DataAddr ? buffer_787 : _GEN_1810; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1812 = 10'h314 == io_BankIO_DataAddr ? buffer_788 : _GEN_1811; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1813 = 10'h315 == io_BankIO_DataAddr ? buffer_789 : _GEN_1812; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1814 = 10'h316 == io_BankIO_DataAddr ? buffer_790 : _GEN_1813; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1815 = 10'h317 == io_BankIO_DataAddr ? buffer_791 : _GEN_1814; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1816 = 10'h318 == io_BankIO_DataAddr ? buffer_792 : _GEN_1815; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1817 = 10'h319 == io_BankIO_DataAddr ? buffer_793 : _GEN_1816; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1818 = 10'h31a == io_BankIO_DataAddr ? buffer_794 : _GEN_1817; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1819 = 10'h31b == io_BankIO_DataAddr ? buffer_795 : _GEN_1818; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1820 = 10'h31c == io_BankIO_DataAddr ? buffer_796 : _GEN_1819; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1821 = 10'h31d == io_BankIO_DataAddr ? buffer_797 : _GEN_1820; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1822 = 10'h31e == io_BankIO_DataAddr ? buffer_798 : _GEN_1821; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1823 = 10'h31f == io_BankIO_DataAddr ? buffer_799 : _GEN_1822; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1824 = 10'h320 == io_BankIO_DataAddr ? buffer_800 : _GEN_1823; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1825 = 10'h321 == io_BankIO_DataAddr ? buffer_801 : _GEN_1824; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1826 = 10'h322 == io_BankIO_DataAddr ? buffer_802 : _GEN_1825; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1827 = 10'h323 == io_BankIO_DataAddr ? buffer_803 : _GEN_1826; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1828 = 10'h324 == io_BankIO_DataAddr ? buffer_804 : _GEN_1827; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1829 = 10'h325 == io_BankIO_DataAddr ? buffer_805 : _GEN_1828; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1830 = 10'h326 == io_BankIO_DataAddr ? buffer_806 : _GEN_1829; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1831 = 10'h327 == io_BankIO_DataAddr ? buffer_807 : _GEN_1830; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1832 = 10'h328 == io_BankIO_DataAddr ? buffer_808 : _GEN_1831; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1833 = 10'h329 == io_BankIO_DataAddr ? buffer_809 : _GEN_1832; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1834 = 10'h32a == io_BankIO_DataAddr ? buffer_810 : _GEN_1833; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1835 = 10'h32b == io_BankIO_DataAddr ? buffer_811 : _GEN_1834; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1836 = 10'h32c == io_BankIO_DataAddr ? buffer_812 : _GEN_1835; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1837 = 10'h32d == io_BankIO_DataAddr ? buffer_813 : _GEN_1836; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1838 = 10'h32e == io_BankIO_DataAddr ? buffer_814 : _GEN_1837; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1839 = 10'h32f == io_BankIO_DataAddr ? buffer_815 : _GEN_1838; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1840 = 10'h330 == io_BankIO_DataAddr ? buffer_816 : _GEN_1839; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1841 = 10'h331 == io_BankIO_DataAddr ? buffer_817 : _GEN_1840; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1842 = 10'h332 == io_BankIO_DataAddr ? buffer_818 : _GEN_1841; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1843 = 10'h333 == io_BankIO_DataAddr ? buffer_819 : _GEN_1842; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1844 = 10'h334 == io_BankIO_DataAddr ? buffer_820 : _GEN_1843; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1845 = 10'h335 == io_BankIO_DataAddr ? buffer_821 : _GEN_1844; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1846 = 10'h336 == io_BankIO_DataAddr ? buffer_822 : _GEN_1845; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1847 = 10'h337 == io_BankIO_DataAddr ? buffer_823 : _GEN_1846; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1848 = 10'h338 == io_BankIO_DataAddr ? buffer_824 : _GEN_1847; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1849 = 10'h339 == io_BankIO_DataAddr ? buffer_825 : _GEN_1848; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1850 = 10'h33a == io_BankIO_DataAddr ? buffer_826 : _GEN_1849; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1851 = 10'h33b == io_BankIO_DataAddr ? buffer_827 : _GEN_1850; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1852 = 10'h33c == io_BankIO_DataAddr ? buffer_828 : _GEN_1851; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1853 = 10'h33d == io_BankIO_DataAddr ? buffer_829 : _GEN_1852; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1854 = 10'h33e == io_BankIO_DataAddr ? buffer_830 : _GEN_1853; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1855 = 10'h33f == io_BankIO_DataAddr ? buffer_831 : _GEN_1854; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1856 = 10'h340 == io_BankIO_DataAddr ? buffer_832 : _GEN_1855; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1857 = 10'h341 == io_BankIO_DataAddr ? buffer_833 : _GEN_1856; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1858 = 10'h342 == io_BankIO_DataAddr ? buffer_834 : _GEN_1857; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1859 = 10'h343 == io_BankIO_DataAddr ? buffer_835 : _GEN_1858; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1860 = 10'h344 == io_BankIO_DataAddr ? buffer_836 : _GEN_1859; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1861 = 10'h345 == io_BankIO_DataAddr ? buffer_837 : _GEN_1860; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1862 = 10'h346 == io_BankIO_DataAddr ? buffer_838 : _GEN_1861; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1863 = 10'h347 == io_BankIO_DataAddr ? buffer_839 : _GEN_1862; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1864 = 10'h348 == io_BankIO_DataAddr ? buffer_840 : _GEN_1863; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1865 = 10'h349 == io_BankIO_DataAddr ? buffer_841 : _GEN_1864; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1866 = 10'h34a == io_BankIO_DataAddr ? buffer_842 : _GEN_1865; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1867 = 10'h34b == io_BankIO_DataAddr ? buffer_843 : _GEN_1866; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1868 = 10'h34c == io_BankIO_DataAddr ? buffer_844 : _GEN_1867; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1869 = 10'h34d == io_BankIO_DataAddr ? buffer_845 : _GEN_1868; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1870 = 10'h34e == io_BankIO_DataAddr ? buffer_846 : _GEN_1869; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1871 = 10'h34f == io_BankIO_DataAddr ? buffer_847 : _GEN_1870; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1872 = 10'h350 == io_BankIO_DataAddr ? buffer_848 : _GEN_1871; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1873 = 10'h351 == io_BankIO_DataAddr ? buffer_849 : _GEN_1872; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1874 = 10'h352 == io_BankIO_DataAddr ? buffer_850 : _GEN_1873; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1875 = 10'h353 == io_BankIO_DataAddr ? buffer_851 : _GEN_1874; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1876 = 10'h354 == io_BankIO_DataAddr ? buffer_852 : _GEN_1875; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1877 = 10'h355 == io_BankIO_DataAddr ? buffer_853 : _GEN_1876; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1878 = 10'h356 == io_BankIO_DataAddr ? buffer_854 : _GEN_1877; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1879 = 10'h357 == io_BankIO_DataAddr ? buffer_855 : _GEN_1878; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1880 = 10'h358 == io_BankIO_DataAddr ? buffer_856 : _GEN_1879; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1881 = 10'h359 == io_BankIO_DataAddr ? buffer_857 : _GEN_1880; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1882 = 10'h35a == io_BankIO_DataAddr ? buffer_858 : _GEN_1881; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1883 = 10'h35b == io_BankIO_DataAddr ? buffer_859 : _GEN_1882; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1884 = 10'h35c == io_BankIO_DataAddr ? buffer_860 : _GEN_1883; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1885 = 10'h35d == io_BankIO_DataAddr ? buffer_861 : _GEN_1884; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1886 = 10'h35e == io_BankIO_DataAddr ? buffer_862 : _GEN_1885; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1887 = 10'h35f == io_BankIO_DataAddr ? buffer_863 : _GEN_1886; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1888 = 10'h360 == io_BankIO_DataAddr ? buffer_864 : _GEN_1887; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1889 = 10'h361 == io_BankIO_DataAddr ? buffer_865 : _GEN_1888; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1890 = 10'h362 == io_BankIO_DataAddr ? buffer_866 : _GEN_1889; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1891 = 10'h363 == io_BankIO_DataAddr ? buffer_867 : _GEN_1890; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1892 = 10'h364 == io_BankIO_DataAddr ? buffer_868 : _GEN_1891; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1893 = 10'h365 == io_BankIO_DataAddr ? buffer_869 : _GEN_1892; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1894 = 10'h366 == io_BankIO_DataAddr ? buffer_870 : _GEN_1893; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1895 = 10'h367 == io_BankIO_DataAddr ? buffer_871 : _GEN_1894; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1896 = 10'h368 == io_BankIO_DataAddr ? buffer_872 : _GEN_1895; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1897 = 10'h369 == io_BankIO_DataAddr ? buffer_873 : _GEN_1896; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1898 = 10'h36a == io_BankIO_DataAddr ? buffer_874 : _GEN_1897; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1899 = 10'h36b == io_BankIO_DataAddr ? buffer_875 : _GEN_1898; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1900 = 10'h36c == io_BankIO_DataAddr ? buffer_876 : _GEN_1899; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1901 = 10'h36d == io_BankIO_DataAddr ? buffer_877 : _GEN_1900; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1902 = 10'h36e == io_BankIO_DataAddr ? buffer_878 : _GEN_1901; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1903 = 10'h36f == io_BankIO_DataAddr ? buffer_879 : _GEN_1902; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1904 = 10'h370 == io_BankIO_DataAddr ? buffer_880 : _GEN_1903; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1905 = 10'h371 == io_BankIO_DataAddr ? buffer_881 : _GEN_1904; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1906 = 10'h372 == io_BankIO_DataAddr ? buffer_882 : _GEN_1905; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1907 = 10'h373 == io_BankIO_DataAddr ? buffer_883 : _GEN_1906; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1908 = 10'h374 == io_BankIO_DataAddr ? buffer_884 : _GEN_1907; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1909 = 10'h375 == io_BankIO_DataAddr ? buffer_885 : _GEN_1908; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1910 = 10'h376 == io_BankIO_DataAddr ? buffer_886 : _GEN_1909; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1911 = 10'h377 == io_BankIO_DataAddr ? buffer_887 : _GEN_1910; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1912 = 10'h378 == io_BankIO_DataAddr ? buffer_888 : _GEN_1911; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1913 = 10'h379 == io_BankIO_DataAddr ? buffer_889 : _GEN_1912; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1914 = 10'h37a == io_BankIO_DataAddr ? buffer_890 : _GEN_1913; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1915 = 10'h37b == io_BankIO_DataAddr ? buffer_891 : _GEN_1914; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1916 = 10'h37c == io_BankIO_DataAddr ? buffer_892 : _GEN_1915; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1917 = 10'h37d == io_BankIO_DataAddr ? buffer_893 : _GEN_1916; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1918 = 10'h37e == io_BankIO_DataAddr ? buffer_894 : _GEN_1917; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1919 = 10'h37f == io_BankIO_DataAddr ? buffer_895 : _GEN_1918; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1920 = 10'h380 == io_BankIO_DataAddr ? buffer_896 : _GEN_1919; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1921 = 10'h381 == io_BankIO_DataAddr ? buffer_897 : _GEN_1920; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1922 = 10'h382 == io_BankIO_DataAddr ? buffer_898 : _GEN_1921; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1923 = 10'h383 == io_BankIO_DataAddr ? buffer_899 : _GEN_1922; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1924 = 10'h384 == io_BankIO_DataAddr ? buffer_900 : _GEN_1923; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1925 = 10'h385 == io_BankIO_DataAddr ? buffer_901 : _GEN_1924; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1926 = 10'h386 == io_BankIO_DataAddr ? buffer_902 : _GEN_1925; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1927 = 10'h387 == io_BankIO_DataAddr ? buffer_903 : _GEN_1926; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1928 = 10'h388 == io_BankIO_DataAddr ? buffer_904 : _GEN_1927; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1929 = 10'h389 == io_BankIO_DataAddr ? buffer_905 : _GEN_1928; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1930 = 10'h38a == io_BankIO_DataAddr ? buffer_906 : _GEN_1929; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1931 = 10'h38b == io_BankIO_DataAddr ? buffer_907 : _GEN_1930; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1932 = 10'h38c == io_BankIO_DataAddr ? buffer_908 : _GEN_1931; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1933 = 10'h38d == io_BankIO_DataAddr ? buffer_909 : _GEN_1932; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1934 = 10'h38e == io_BankIO_DataAddr ? buffer_910 : _GEN_1933; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1935 = 10'h38f == io_BankIO_DataAddr ? buffer_911 : _GEN_1934; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1936 = 10'h390 == io_BankIO_DataAddr ? buffer_912 : _GEN_1935; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1937 = 10'h391 == io_BankIO_DataAddr ? buffer_913 : _GEN_1936; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1938 = 10'h392 == io_BankIO_DataAddr ? buffer_914 : _GEN_1937; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1939 = 10'h393 == io_BankIO_DataAddr ? buffer_915 : _GEN_1938; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1940 = 10'h394 == io_BankIO_DataAddr ? buffer_916 : _GEN_1939; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1941 = 10'h395 == io_BankIO_DataAddr ? buffer_917 : _GEN_1940; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1942 = 10'h396 == io_BankIO_DataAddr ? buffer_918 : _GEN_1941; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1943 = 10'h397 == io_BankIO_DataAddr ? buffer_919 : _GEN_1942; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1944 = 10'h398 == io_BankIO_DataAddr ? buffer_920 : _GEN_1943; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1945 = 10'h399 == io_BankIO_DataAddr ? buffer_921 : _GEN_1944; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1946 = 10'h39a == io_BankIO_DataAddr ? buffer_922 : _GEN_1945; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1947 = 10'h39b == io_BankIO_DataAddr ? buffer_923 : _GEN_1946; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1948 = 10'h39c == io_BankIO_DataAddr ? buffer_924 : _GEN_1947; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1949 = 10'h39d == io_BankIO_DataAddr ? buffer_925 : _GEN_1948; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1950 = 10'h39e == io_BankIO_DataAddr ? buffer_926 : _GEN_1949; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1951 = 10'h39f == io_BankIO_DataAddr ? buffer_927 : _GEN_1950; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1952 = 10'h3a0 == io_BankIO_DataAddr ? buffer_928 : _GEN_1951; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1953 = 10'h3a1 == io_BankIO_DataAddr ? buffer_929 : _GEN_1952; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1954 = 10'h3a2 == io_BankIO_DataAddr ? buffer_930 : _GEN_1953; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1955 = 10'h3a3 == io_BankIO_DataAddr ? buffer_931 : _GEN_1954; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1956 = 10'h3a4 == io_BankIO_DataAddr ? buffer_932 : _GEN_1955; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1957 = 10'h3a5 == io_BankIO_DataAddr ? buffer_933 : _GEN_1956; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1958 = 10'h3a6 == io_BankIO_DataAddr ? buffer_934 : _GEN_1957; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1959 = 10'h3a7 == io_BankIO_DataAddr ? buffer_935 : _GEN_1958; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1960 = 10'h3a8 == io_BankIO_DataAddr ? buffer_936 : _GEN_1959; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1961 = 10'h3a9 == io_BankIO_DataAddr ? buffer_937 : _GEN_1960; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1962 = 10'h3aa == io_BankIO_DataAddr ? buffer_938 : _GEN_1961; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1963 = 10'h3ab == io_BankIO_DataAddr ? buffer_939 : _GEN_1962; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1964 = 10'h3ac == io_BankIO_DataAddr ? buffer_940 : _GEN_1963; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1965 = 10'h3ad == io_BankIO_DataAddr ? buffer_941 : _GEN_1964; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1966 = 10'h3ae == io_BankIO_DataAddr ? buffer_942 : _GEN_1965; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1967 = 10'h3af == io_BankIO_DataAddr ? buffer_943 : _GEN_1966; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1968 = 10'h3b0 == io_BankIO_DataAddr ? buffer_944 : _GEN_1967; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1969 = 10'h3b1 == io_BankIO_DataAddr ? buffer_945 : _GEN_1968; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1970 = 10'h3b2 == io_BankIO_DataAddr ? buffer_946 : _GEN_1969; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1971 = 10'h3b3 == io_BankIO_DataAddr ? buffer_947 : _GEN_1970; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1972 = 10'h3b4 == io_BankIO_DataAddr ? buffer_948 : _GEN_1971; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1973 = 10'h3b5 == io_BankIO_DataAddr ? buffer_949 : _GEN_1972; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1974 = 10'h3b6 == io_BankIO_DataAddr ? buffer_950 : _GEN_1973; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1975 = 10'h3b7 == io_BankIO_DataAddr ? buffer_951 : _GEN_1974; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1976 = 10'h3b8 == io_BankIO_DataAddr ? buffer_952 : _GEN_1975; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1977 = 10'h3b9 == io_BankIO_DataAddr ? buffer_953 : _GEN_1976; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1978 = 10'h3ba == io_BankIO_DataAddr ? buffer_954 : _GEN_1977; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1979 = 10'h3bb == io_BankIO_DataAddr ? buffer_955 : _GEN_1978; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1980 = 10'h3bc == io_BankIO_DataAddr ? buffer_956 : _GEN_1979; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1981 = 10'h3bd == io_BankIO_DataAddr ? buffer_957 : _GEN_1980; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1982 = 10'h3be == io_BankIO_DataAddr ? buffer_958 : _GEN_1981; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1983 = 10'h3bf == io_BankIO_DataAddr ? buffer_959 : _GEN_1982; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1984 = 10'h3c0 == io_BankIO_DataAddr ? buffer_960 : _GEN_1983; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1985 = 10'h3c1 == io_BankIO_DataAddr ? buffer_961 : _GEN_1984; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1986 = 10'h3c2 == io_BankIO_DataAddr ? buffer_962 : _GEN_1985; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1987 = 10'h3c3 == io_BankIO_DataAddr ? buffer_963 : _GEN_1986; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1988 = 10'h3c4 == io_BankIO_DataAddr ? buffer_964 : _GEN_1987; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1989 = 10'h3c5 == io_BankIO_DataAddr ? buffer_965 : _GEN_1988; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1990 = 10'h3c6 == io_BankIO_DataAddr ? buffer_966 : _GEN_1989; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1991 = 10'h3c7 == io_BankIO_DataAddr ? buffer_967 : _GEN_1990; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1992 = 10'h3c8 == io_BankIO_DataAddr ? buffer_968 : _GEN_1991; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1993 = 10'h3c9 == io_BankIO_DataAddr ? buffer_969 : _GEN_1992; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1994 = 10'h3ca == io_BankIO_DataAddr ? buffer_970 : _GEN_1993; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1995 = 10'h3cb == io_BankIO_DataAddr ? buffer_971 : _GEN_1994; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1996 = 10'h3cc == io_BankIO_DataAddr ? buffer_972 : _GEN_1995; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1997 = 10'h3cd == io_BankIO_DataAddr ? buffer_973 : _GEN_1996; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1998 = 10'h3ce == io_BankIO_DataAddr ? buffer_974 : _GEN_1997; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_1999 = 10'h3cf == io_BankIO_DataAddr ? buffer_975 : _GEN_1998; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2000 = 10'h3d0 == io_BankIO_DataAddr ? buffer_976 : _GEN_1999; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2001 = 10'h3d1 == io_BankIO_DataAddr ? buffer_977 : _GEN_2000; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2002 = 10'h3d2 == io_BankIO_DataAddr ? buffer_978 : _GEN_2001; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2003 = 10'h3d3 == io_BankIO_DataAddr ? buffer_979 : _GEN_2002; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2004 = 10'h3d4 == io_BankIO_DataAddr ? buffer_980 : _GEN_2003; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2005 = 10'h3d5 == io_BankIO_DataAddr ? buffer_981 : _GEN_2004; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2006 = 10'h3d6 == io_BankIO_DataAddr ? buffer_982 : _GEN_2005; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2007 = 10'h3d7 == io_BankIO_DataAddr ? buffer_983 : _GEN_2006; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2008 = 10'h3d8 == io_BankIO_DataAddr ? buffer_984 : _GEN_2007; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2009 = 10'h3d9 == io_BankIO_DataAddr ? buffer_985 : _GEN_2008; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2010 = 10'h3da == io_BankIO_DataAddr ? buffer_986 : _GEN_2009; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2011 = 10'h3db == io_BankIO_DataAddr ? buffer_987 : _GEN_2010; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2012 = 10'h3dc == io_BankIO_DataAddr ? buffer_988 : _GEN_2011; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2013 = 10'h3dd == io_BankIO_DataAddr ? buffer_989 : _GEN_2012; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2014 = 10'h3de == io_BankIO_DataAddr ? buffer_990 : _GEN_2013; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2015 = 10'h3df == io_BankIO_DataAddr ? buffer_991 : _GEN_2014; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2016 = 10'h3e0 == io_BankIO_DataAddr ? buffer_992 : _GEN_2015; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2017 = 10'h3e1 == io_BankIO_DataAddr ? buffer_993 : _GEN_2016; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2018 = 10'h3e2 == io_BankIO_DataAddr ? buffer_994 : _GEN_2017; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2019 = 10'h3e3 == io_BankIO_DataAddr ? buffer_995 : _GEN_2018; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2020 = 10'h3e4 == io_BankIO_DataAddr ? buffer_996 : _GEN_2019; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2021 = 10'h3e5 == io_BankIO_DataAddr ? buffer_997 : _GEN_2020; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2022 = 10'h3e6 == io_BankIO_DataAddr ? buffer_998 : _GEN_2021; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2023 = 10'h3e7 == io_BankIO_DataAddr ? buffer_999 : _GEN_2022; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2024 = 10'h3e8 == io_BankIO_DataAddr ? buffer_1000 : _GEN_2023; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2025 = 10'h3e9 == io_BankIO_DataAddr ? buffer_1001 : _GEN_2024; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2026 = 10'h3ea == io_BankIO_DataAddr ? buffer_1002 : _GEN_2025; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2027 = 10'h3eb == io_BankIO_DataAddr ? buffer_1003 : _GEN_2026; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2028 = 10'h3ec == io_BankIO_DataAddr ? buffer_1004 : _GEN_2027; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2029 = 10'h3ed == io_BankIO_DataAddr ? buffer_1005 : _GEN_2028; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2030 = 10'h3ee == io_BankIO_DataAddr ? buffer_1006 : _GEN_2029; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2031 = 10'h3ef == io_BankIO_DataAddr ? buffer_1007 : _GEN_2030; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2032 = 10'h3f0 == io_BankIO_DataAddr ? buffer_1008 : _GEN_2031; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2033 = 10'h3f1 == io_BankIO_DataAddr ? buffer_1009 : _GEN_2032; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2034 = 10'h3f2 == io_BankIO_DataAddr ? buffer_1010 : _GEN_2033; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2035 = 10'h3f3 == io_BankIO_DataAddr ? buffer_1011 : _GEN_2034; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2036 = 10'h3f4 == io_BankIO_DataAddr ? buffer_1012 : _GEN_2035; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2037 = 10'h3f5 == io_BankIO_DataAddr ? buffer_1013 : _GEN_2036; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2038 = 10'h3f6 == io_BankIO_DataAddr ? buffer_1014 : _GEN_2037; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2039 = 10'h3f7 == io_BankIO_DataAddr ? buffer_1015 : _GEN_2038; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2040 = 10'h3f8 == io_BankIO_DataAddr ? buffer_1016 : _GEN_2039; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2041 = 10'h3f9 == io_BankIO_DataAddr ? buffer_1017 : _GEN_2040; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2042 = 10'h3fa == io_BankIO_DataAddr ? buffer_1018 : _GEN_2041; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2043 = 10'h3fb == io_BankIO_DataAddr ? buffer_1019 : _GEN_2042; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2044 = 10'h3fc == io_BankIO_DataAddr ? buffer_1020 : _GEN_2043; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2045 = 10'h3fd == io_BankIO_DataAddr ? buffer_1021 : _GEN_2044; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2046 = 10'h3fe == io_BankIO_DataAddr ? buffer_1022 : _GEN_2045; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_2047 = 10'h3ff == io_BankIO_DataAddr ? buffer_1023 : _GEN_2046; // @[OuterBuffer.scala 27:{25,25}]
  wire [15:0] _GEN_3072 = ~io_BankIO_ReadWrite ? 16'h0 : _GEN_2047; // @[OuterBuffer.scala 22:21 24:43 27:25]
  assign io_BankIO_DataOut = io_BankIO_Enable ? _GEN_3072 : 16'h0; // @[OuterBuffer.scala 22:21 23:37]
  always @(posedge clock) begin
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_0 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_0 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_2 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_2 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_3 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_3 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_4 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_4 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_5 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_5 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_6 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_6 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_7 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_7 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_8 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_8 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_9 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_9 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_10 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_10 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_11 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_11 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_12 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_12 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_13 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_13 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_14 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_14 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_15 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_15 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_16 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h10 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_16 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_17 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h11 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_17 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_18 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h12 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_18 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_19 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h13 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_19 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_20 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h14 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_20 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_21 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h15 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_21 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_22 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h16 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_22 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_23 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h17 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_23 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_24 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h18 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_24 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_25 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h19 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_25 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_26 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_26 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_27 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_27 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_28 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_28 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_29 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_29 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_30 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_30 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_31 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_31 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_32 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h20 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_32 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_33 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h21 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_33 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_34 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h22 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_34 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_35 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h23 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_35 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_36 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h24 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_36 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_37 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h25 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_37 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_38 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h26 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_38 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_39 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h27 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_39 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_40 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h28 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_40 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_41 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h29 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_41 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_42 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_42 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_43 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_43 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_44 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_44 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_45 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_45 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_46 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_46 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_47 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_47 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_48 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h30 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_48 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_49 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h31 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_49 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_50 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h32 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_50 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_51 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h33 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_51 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_52 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h34 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_52 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_53 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h35 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_53 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_54 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h36 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_54 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_55 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h37 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_55 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_56 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h38 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_56 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_57 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h39 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_57 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_58 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_58 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_59 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_59 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_60 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_60 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_61 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_61 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_62 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_62 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_63 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_63 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_64 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h40 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_64 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_65 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h41 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_65 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_66 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h42 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_66 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_67 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h43 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_67 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_68 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h44 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_68 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_69 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h45 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_69 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_70 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h46 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_70 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_71 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h47 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_71 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_72 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h48 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_72 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_73 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h49 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_73 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_74 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h4a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_74 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_75 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h4b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_75 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_76 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h4c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_76 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_77 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h4d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_77 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_78 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h4e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_78 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_79 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h4f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_79 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_80 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h50 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_80 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_81 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h51 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_81 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_82 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h52 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_82 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_83 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h53 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_83 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_84 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h54 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_84 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_85 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h55 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_85 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_86 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h56 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_86 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_87 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h57 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_87 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_88 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h58 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_88 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_89 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h59 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_89 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_90 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h5a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_90 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_91 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h5b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_91 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_92 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h5c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_92 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_93 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h5d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_93 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_94 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h5e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_94 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_95 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h5f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_95 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_96 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h60 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_96 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_97 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h61 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_97 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_98 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h62 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_98 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_99 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h63 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_99 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_100 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h64 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_100 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_101 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h65 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_101 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_102 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h66 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_102 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_103 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h67 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_103 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_104 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h68 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_104 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_105 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h69 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_105 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_106 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h6a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_106 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_107 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h6b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_107 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_108 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h6c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_108 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_109 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h6d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_109 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_110 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h6e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_110 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_111 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h6f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_111 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_112 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h70 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_112 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_113 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h71 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_113 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_114 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h72 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_114 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_115 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h73 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_115 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_116 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h74 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_116 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_117 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h75 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_117 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_118 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h76 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_118 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_119 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h77 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_119 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_120 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h78 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_120 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_121 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h79 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_121 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_122 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h7a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_122 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_123 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h7b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_123 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_124 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h7c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_124 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_125 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h7d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_125 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_126 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h7e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_126 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_127 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h7f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_127 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_128 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h80 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_128 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_129 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h81 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_129 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_130 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h82 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_130 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_131 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h83 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_131 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_132 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h84 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_132 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_133 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h85 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_133 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_134 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h86 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_134 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_135 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h87 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_135 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_136 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h88 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_136 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_137 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h89 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_137 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_138 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h8a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_138 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_139 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h8b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_139 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_140 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h8c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_140 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_141 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h8d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_141 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_142 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h8e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_142 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_143 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h8f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_143 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_144 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h90 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_144 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_145 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h91 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_145 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_146 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h92 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_146 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_147 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h93 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_147 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_148 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h94 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_148 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_149 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h95 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_149 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_150 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h96 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_150 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_151 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h97 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_151 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_152 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h98 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_152 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_153 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h99 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_153 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_154 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h9a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_154 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_155 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h9b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_155 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_156 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h9c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_156 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_157 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h9d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_157 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_158 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h9e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_158 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_159 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h9f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_159 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_160 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_160 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_161 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_161 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_162 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_162 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_163 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_163 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_164 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_164 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_165 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_165 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_166 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_166 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_167 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_167 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_168 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_168 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_169 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'ha9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_169 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_170 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'haa == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_170 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_171 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hab == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_171 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_172 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hac == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_172 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_173 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'had == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_173 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_174 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hae == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_174 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_175 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'haf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_175 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_176 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_176 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_177 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_177 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_178 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_178 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_179 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_179 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_180 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_180 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_181 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_181 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_182 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_182 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_183 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_183 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_184 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_184 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_185 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hb9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_185 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_186 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hba == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_186 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_187 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hbb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_187 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_188 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hbc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_188 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_189 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hbd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_189 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_190 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hbe == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_190 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_191 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hbf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_191 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_192 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_192 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_193 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_193 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_194 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_194 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_195 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_195 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_196 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_196 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_197 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_197 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_198 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_198 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_199 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_199 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_200 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_200 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_201 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hc9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_201 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_202 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hca == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_202 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_203 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hcb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_203 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_204 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hcc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_204 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_205 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hcd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_205 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_206 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hce == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_206 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_207 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hcf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_207 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_208 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_208 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_209 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_209 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_210 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_210 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_211 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_211 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_212 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_212 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_213 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_213 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_214 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_214 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_215 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_215 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_216 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_216 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_217 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hd9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_217 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_218 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hda == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_218 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_219 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hdb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_219 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_220 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hdc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_220 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_221 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hdd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_221 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_222 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hde == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_222 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_223 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hdf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_223 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_224 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_224 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_225 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_225 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_226 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_226 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_227 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_227 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_228 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_228 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_229 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_229 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_230 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_230 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_231 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_231 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_232 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_232 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_233 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'he9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_233 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_234 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hea == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_234 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_235 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'heb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_235 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_236 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hec == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_236 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_237 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hed == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_237 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_238 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hee == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_238 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_239 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hef == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_239 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_240 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_240 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_241 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_241 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_242 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_242 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_243 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_243 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_244 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_244 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_245 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_245 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_246 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_246 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_247 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_247 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_248 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_248 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_249 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hf9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_249 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_250 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hfa == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_250 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_251 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hfb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_251 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_252 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hfc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_252 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_253 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hfd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_253 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_254 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hfe == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_254 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_255 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'hff == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_255 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_256 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h100 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_256 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_257 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h101 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_257 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_258 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h102 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_258 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_259 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h103 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_259 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_260 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h104 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_260 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_261 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h105 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_261 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_262 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h106 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_262 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_263 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h107 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_263 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_264 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h108 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_264 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_265 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h109 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_265 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_266 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h10a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_266 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_267 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h10b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_267 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_268 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h10c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_268 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_269 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h10d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_269 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_270 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h10e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_270 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_271 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h10f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_271 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_272 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h110 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_272 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_273 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h111 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_273 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_274 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h112 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_274 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_275 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h113 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_275 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_276 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h114 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_276 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_277 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h115 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_277 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_278 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h116 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_278 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_279 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h117 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_279 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_280 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h118 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_280 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_281 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h119 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_281 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_282 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h11a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_282 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_283 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h11b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_283 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_284 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h11c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_284 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_285 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h11d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_285 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_286 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h11e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_286 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_287 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h11f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_287 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_288 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h120 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_288 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_289 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h121 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_289 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_290 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h122 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_290 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_291 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h123 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_291 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_292 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h124 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_292 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_293 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h125 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_293 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_294 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h126 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_294 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_295 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h127 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_295 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_296 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h128 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_296 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_297 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h129 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_297 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_298 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h12a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_298 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_299 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h12b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_299 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_300 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h12c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_300 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_301 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h12d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_301 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_302 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h12e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_302 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_303 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h12f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_303 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_304 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h130 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_304 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_305 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h131 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_305 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_306 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h132 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_306 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_307 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h133 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_307 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_308 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h134 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_308 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_309 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h135 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_309 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_310 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h136 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_310 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_311 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h137 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_311 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_312 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h138 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_312 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_313 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h139 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_313 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_314 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h13a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_314 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_315 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h13b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_315 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_316 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h13c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_316 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_317 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h13d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_317 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_318 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h13e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_318 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_319 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h13f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_319 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_320 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h140 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_320 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_321 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h141 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_321 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_322 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h142 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_322 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_323 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h143 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_323 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_324 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h144 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_324 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_325 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h145 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_325 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_326 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h146 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_326 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_327 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h147 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_327 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_328 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h148 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_328 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_329 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h149 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_329 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_330 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h14a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_330 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_331 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h14b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_331 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_332 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h14c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_332 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_333 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h14d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_333 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_334 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h14e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_334 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_335 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h14f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_335 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_336 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h150 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_336 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_337 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h151 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_337 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_338 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h152 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_338 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_339 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h153 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_339 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_340 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h154 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_340 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_341 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h155 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_341 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_342 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h156 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_342 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_343 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h157 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_343 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_344 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h158 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_344 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_345 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h159 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_345 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_346 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h15a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_346 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_347 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h15b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_347 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_348 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h15c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_348 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_349 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h15d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_349 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_350 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h15e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_350 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_351 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h15f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_351 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_352 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h160 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_352 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_353 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h161 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_353 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_354 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h162 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_354 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_355 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h163 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_355 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_356 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h164 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_356 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_357 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h165 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_357 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_358 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h166 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_358 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_359 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h167 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_359 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_360 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h168 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_360 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_361 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h169 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_361 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_362 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h16a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_362 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_363 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h16b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_363 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_364 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h16c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_364 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_365 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h16d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_365 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_366 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h16e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_366 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_367 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h16f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_367 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_368 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h170 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_368 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_369 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h171 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_369 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_370 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h172 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_370 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_371 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h173 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_371 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_372 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h174 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_372 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_373 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h175 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_373 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_374 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h176 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_374 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_375 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h177 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_375 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_376 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h178 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_376 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_377 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h179 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_377 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_378 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h17a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_378 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_379 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h17b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_379 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_380 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h17c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_380 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_381 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h17d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_381 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_382 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h17e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_382 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_383 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h17f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_383 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_384 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h180 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_384 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_385 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h181 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_385 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_386 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h182 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_386 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_387 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h183 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_387 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_388 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h184 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_388 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_389 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h185 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_389 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_390 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h186 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_390 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_391 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h187 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_391 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_392 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h188 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_392 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_393 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h189 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_393 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_394 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h18a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_394 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_395 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h18b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_395 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_396 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h18c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_396 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_397 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h18d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_397 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_398 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h18e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_398 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_399 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h18f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_399 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_400 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h190 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_400 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_401 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h191 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_401 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_402 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h192 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_402 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_403 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h193 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_403 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_404 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h194 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_404 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_405 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h195 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_405 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_406 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h196 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_406 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_407 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h197 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_407 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_408 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h198 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_408 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_409 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h199 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_409 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_410 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h19a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_410 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_411 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h19b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_411 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_412 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h19c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_412 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_413 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h19d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_413 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_414 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h19e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_414 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_415 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h19f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_415 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_416 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_416 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_417 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_417 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_418 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_418 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_419 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_419 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_420 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_420 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_421 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_421 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_422 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_422 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_423 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_423 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_424 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_424 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_425 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1a9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_425 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_426 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1aa == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_426 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_427 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ab == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_427 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_428 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ac == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_428 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_429 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ad == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_429 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_430 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ae == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_430 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_431 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1af == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_431 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_432 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_432 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_433 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_433 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_434 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_434 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_435 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_435 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_436 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_436 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_437 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_437 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_438 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_438 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_439 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_439 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_440 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_440 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_441 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1b9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_441 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_442 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ba == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_442 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_443 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1bb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_443 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_444 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1bc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_444 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_445 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1bd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_445 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_446 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1be == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_446 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_447 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1bf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_447 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_448 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_448 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_449 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_449 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_450 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_450 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_451 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_451 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_452 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_452 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_453 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_453 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_454 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_454 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_455 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_455 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_456 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_456 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_457 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1c9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_457 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_458 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ca == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_458 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_459 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1cb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_459 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_460 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1cc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_460 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_461 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1cd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_461 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_462 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ce == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_462 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_463 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1cf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_463 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_464 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_464 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_465 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_465 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_466 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_466 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_467 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_467 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_468 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_468 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_469 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_469 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_470 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_470 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_471 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_471 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_472 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_472 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_473 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1d9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_473 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_474 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1da == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_474 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_475 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1db == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_475 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_476 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1dc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_476 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_477 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1dd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_477 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_478 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1de == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_478 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_479 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1df == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_479 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_480 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_480 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_481 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_481 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_482 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_482 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_483 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_483 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_484 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_484 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_485 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_485 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_486 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_486 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_487 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_487 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_488 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_488 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_489 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1e9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_489 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_490 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ea == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_490 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_491 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1eb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_491 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_492 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ec == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_492 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_493 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ed == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_493 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_494 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ee == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_494 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_495 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ef == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_495 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_496 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_496 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_497 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_497 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_498 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_498 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_499 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_499 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_500 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_500 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_501 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_501 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_502 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_502 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_503 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_503 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_504 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_504 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_505 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1f9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_505 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_506 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1fa == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_506 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_507 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1fb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_507 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_508 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1fc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_508 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_509 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1fd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_509 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_510 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1fe == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_510 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_511 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h1ff == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_511 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_512 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h200 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_512 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_513 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h201 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_513 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_514 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h202 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_514 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_515 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h203 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_515 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_516 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h204 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_516 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_517 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h205 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_517 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_518 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h206 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_518 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_519 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h207 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_519 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_520 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h208 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_520 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_521 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h209 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_521 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_522 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h20a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_522 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_523 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h20b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_523 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_524 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h20c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_524 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_525 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h20d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_525 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_526 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h20e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_526 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_527 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h20f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_527 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_528 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h210 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_528 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_529 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h211 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_529 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_530 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h212 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_530 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_531 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h213 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_531 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_532 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h214 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_532 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_533 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h215 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_533 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_534 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h216 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_534 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_535 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h217 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_535 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_536 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h218 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_536 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_537 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h219 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_537 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_538 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h21a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_538 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_539 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h21b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_539 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_540 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h21c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_540 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_541 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h21d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_541 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_542 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h21e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_542 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_543 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h21f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_543 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_544 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h220 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_544 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_545 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h221 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_545 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_546 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h222 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_546 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_547 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h223 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_547 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_548 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h224 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_548 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_549 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h225 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_549 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_550 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h226 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_550 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_551 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h227 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_551 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_552 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h228 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_552 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_553 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h229 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_553 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_554 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h22a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_554 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_555 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h22b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_555 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_556 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h22c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_556 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_557 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h22d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_557 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_558 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h22e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_558 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_559 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h22f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_559 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_560 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h230 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_560 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_561 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h231 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_561 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_562 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h232 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_562 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_563 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h233 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_563 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_564 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h234 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_564 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_565 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h235 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_565 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_566 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h236 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_566 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_567 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h237 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_567 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_568 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h238 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_568 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_569 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h239 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_569 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_570 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h23a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_570 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_571 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h23b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_571 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_572 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h23c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_572 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_573 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h23d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_573 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_574 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h23e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_574 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_575 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h23f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_575 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_576 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h240 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_576 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_577 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h241 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_577 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_578 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h242 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_578 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_579 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h243 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_579 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_580 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h244 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_580 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_581 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h245 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_581 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_582 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h246 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_582 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_583 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h247 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_583 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_584 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h248 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_584 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_585 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h249 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_585 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_586 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h24a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_586 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_587 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h24b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_587 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_588 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h24c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_588 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_589 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h24d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_589 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_590 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h24e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_590 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_591 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h24f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_591 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_592 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h250 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_592 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_593 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h251 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_593 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_594 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h252 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_594 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_595 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h253 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_595 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_596 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h254 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_596 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_597 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h255 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_597 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_598 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h256 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_598 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_599 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h257 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_599 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_600 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h258 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_600 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_601 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h259 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_601 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_602 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h25a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_602 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_603 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h25b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_603 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_604 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h25c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_604 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_605 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h25d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_605 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_606 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h25e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_606 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_607 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h25f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_607 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_608 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h260 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_608 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_609 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h261 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_609 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_610 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h262 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_610 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_611 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h263 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_611 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_612 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h264 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_612 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_613 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h265 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_613 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_614 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h266 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_614 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_615 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h267 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_615 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_616 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h268 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_616 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_617 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h269 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_617 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_618 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h26a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_618 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_619 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h26b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_619 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_620 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h26c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_620 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_621 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h26d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_621 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_622 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h26e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_622 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_623 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h26f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_623 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_624 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h270 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_624 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_625 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h271 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_625 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_626 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h272 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_626 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_627 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h273 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_627 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_628 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h274 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_628 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_629 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h275 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_629 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_630 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h276 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_630 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_631 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h277 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_631 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_632 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h278 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_632 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_633 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h279 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_633 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_634 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h27a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_634 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_635 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h27b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_635 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_636 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h27c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_636 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_637 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h27d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_637 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_638 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h27e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_638 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_639 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h27f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_639 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_640 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h280 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_640 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_641 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h281 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_641 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_642 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h282 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_642 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_643 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h283 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_643 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_644 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h284 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_644 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_645 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h285 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_645 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_646 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h286 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_646 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_647 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h287 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_647 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_648 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h288 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_648 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_649 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h289 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_649 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_650 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h28a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_650 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_651 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h28b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_651 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_652 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h28c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_652 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_653 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h28d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_653 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_654 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h28e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_654 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_655 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h28f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_655 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_656 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h290 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_656 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_657 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h291 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_657 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_658 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h292 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_658 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_659 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h293 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_659 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_660 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h294 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_660 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_661 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h295 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_661 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_662 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h296 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_662 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_663 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h297 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_663 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_664 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h298 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_664 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_665 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h299 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_665 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_666 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h29a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_666 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_667 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h29b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_667 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_668 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h29c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_668 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_669 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h29d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_669 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_670 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h29e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_670 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_671 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h29f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_671 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_672 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_672 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_673 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_673 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_674 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_674 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_675 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_675 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_676 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_676 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_677 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_677 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_678 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_678 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_679 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_679 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_680 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_680 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_681 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2a9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_681 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_682 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2aa == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_682 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_683 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ab == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_683 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_684 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ac == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_684 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_685 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ad == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_685 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_686 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ae == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_686 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_687 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2af == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_687 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_688 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_688 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_689 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_689 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_690 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_690 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_691 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_691 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_692 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_692 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_693 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_693 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_694 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_694 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_695 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_695 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_696 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_696 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_697 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2b9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_697 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_698 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ba == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_698 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_699 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2bb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_699 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_700 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2bc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_700 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_701 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2bd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_701 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_702 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2be == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_702 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_703 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2bf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_703 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_704 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_704 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_705 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_705 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_706 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_706 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_707 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_707 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_708 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_708 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_709 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_709 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_710 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_710 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_711 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_711 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_712 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_712 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_713 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2c9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_713 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_714 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ca == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_714 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_715 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2cb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_715 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_716 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2cc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_716 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_717 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2cd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_717 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_718 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ce == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_718 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_719 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2cf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_719 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_720 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_720 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_721 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_721 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_722 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_722 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_723 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_723 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_724 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_724 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_725 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_725 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_726 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_726 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_727 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_727 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_728 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_728 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_729 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2d9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_729 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_730 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2da == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_730 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_731 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2db == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_731 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_732 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2dc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_732 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_733 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2dd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_733 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_734 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2de == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_734 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_735 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2df == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_735 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_736 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_736 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_737 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_737 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_738 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_738 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_739 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_739 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_740 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_740 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_741 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_741 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_742 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_742 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_743 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_743 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_744 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_744 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_745 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2e9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_745 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_746 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ea == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_746 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_747 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2eb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_747 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_748 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ec == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_748 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_749 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ed == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_749 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_750 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ee == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_750 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_751 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ef == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_751 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_752 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_752 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_753 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_753 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_754 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_754 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_755 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_755 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_756 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_756 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_757 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_757 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_758 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_758 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_759 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_759 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_760 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_760 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_761 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2f9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_761 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_762 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2fa == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_762 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_763 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2fb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_763 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_764 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2fc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_764 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_765 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2fd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_765 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_766 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2fe == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_766 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_767 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h2ff == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_767 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_768 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h300 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_768 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_769 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h301 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_769 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_770 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h302 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_770 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_771 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h303 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_771 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_772 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h304 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_772 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_773 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h305 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_773 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_774 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h306 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_774 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_775 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h307 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_775 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_776 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h308 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_776 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_777 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h309 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_777 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_778 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h30a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_778 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_779 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h30b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_779 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_780 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h30c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_780 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_781 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h30d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_781 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_782 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h30e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_782 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_783 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h30f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_783 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_784 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h310 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_784 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_785 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h311 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_785 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_786 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h312 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_786 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_787 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h313 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_787 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_788 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h314 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_788 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_789 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h315 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_789 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_790 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h316 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_790 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_791 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h317 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_791 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_792 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h318 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_792 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_793 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h319 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_793 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_794 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h31a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_794 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_795 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h31b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_795 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_796 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h31c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_796 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_797 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h31d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_797 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_798 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h31e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_798 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_799 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h31f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_799 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_800 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h320 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_800 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_801 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h321 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_801 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_802 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h322 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_802 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_803 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h323 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_803 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_804 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h324 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_804 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_805 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h325 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_805 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_806 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h326 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_806 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_807 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h327 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_807 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_808 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h328 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_808 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_809 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h329 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_809 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_810 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h32a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_810 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_811 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h32b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_811 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_812 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h32c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_812 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_813 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h32d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_813 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_814 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h32e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_814 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_815 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h32f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_815 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_816 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h330 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_816 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_817 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h331 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_817 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_818 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h332 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_818 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_819 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h333 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_819 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_820 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h334 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_820 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_821 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h335 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_821 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_822 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h336 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_822 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_823 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h337 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_823 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_824 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h338 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_824 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_825 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h339 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_825 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_826 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h33a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_826 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_827 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h33b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_827 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_828 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h33c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_828 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_829 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h33d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_829 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_830 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h33e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_830 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_831 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h33f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_831 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_832 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h340 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_832 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_833 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h341 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_833 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_834 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h342 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_834 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_835 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h343 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_835 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_836 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h344 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_836 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_837 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h345 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_837 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_838 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h346 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_838 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_839 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h347 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_839 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_840 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h348 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_840 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_841 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h349 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_841 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_842 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h34a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_842 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_843 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h34b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_843 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_844 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h34c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_844 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_845 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h34d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_845 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_846 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h34e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_846 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_847 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h34f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_847 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_848 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h350 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_848 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_849 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h351 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_849 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_850 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h352 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_850 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_851 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h353 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_851 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_852 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h354 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_852 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_853 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h355 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_853 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_854 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h356 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_854 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_855 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h357 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_855 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_856 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h358 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_856 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_857 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h359 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_857 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_858 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h35a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_858 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_859 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h35b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_859 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_860 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h35c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_860 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_861 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h35d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_861 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_862 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h35e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_862 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_863 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h35f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_863 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_864 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h360 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_864 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_865 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h361 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_865 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_866 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h362 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_866 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_867 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h363 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_867 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_868 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h364 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_868 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_869 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h365 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_869 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_870 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h366 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_870 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_871 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h367 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_871 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_872 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h368 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_872 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_873 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h369 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_873 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_874 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h36a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_874 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_875 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h36b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_875 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_876 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h36c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_876 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_877 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h36d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_877 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_878 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h36e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_878 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_879 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h36f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_879 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_880 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h370 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_880 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_881 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h371 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_881 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_882 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h372 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_882 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_883 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h373 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_883 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_884 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h374 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_884 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_885 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h375 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_885 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_886 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h376 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_886 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_887 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h377 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_887 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_888 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h378 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_888 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_889 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h379 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_889 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_890 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h37a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_890 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_891 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h37b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_891 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_892 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h37c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_892 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_893 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h37d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_893 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_894 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h37e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_894 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_895 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h37f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_895 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_896 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h380 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_896 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_897 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h381 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_897 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_898 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h382 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_898 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_899 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h383 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_899 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_900 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h384 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_900 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_901 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h385 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_901 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_902 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h386 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_902 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_903 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h387 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_903 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_904 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h388 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_904 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_905 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h389 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_905 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_906 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h38a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_906 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_907 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h38b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_907 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_908 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h38c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_908 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_909 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h38d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_909 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_910 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h38e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_910 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_911 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h38f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_911 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_912 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h390 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_912 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_913 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h391 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_913 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_914 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h392 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_914 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_915 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h393 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_915 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_916 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h394 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_916 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_917 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h395 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_917 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_918 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h396 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_918 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_919 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h397 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_919 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_920 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h398 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_920 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_921 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h399 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_921 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_922 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h39a == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_922 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_923 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h39b == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_923 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_924 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h39c == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_924 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_925 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h39d == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_925 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_926 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h39e == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_926 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_927 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h39f == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_927 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_928 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_928 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_929 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_929 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_930 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_930 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_931 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_931 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_932 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_932 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_933 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_933 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_934 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_934 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_935 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_935 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_936 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_936 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_937 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3a9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_937 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_938 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3aa == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_938 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_939 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ab == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_939 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_940 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ac == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_940 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_941 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ad == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_941 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_942 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ae == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_942 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_943 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3af == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_943 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_944 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_944 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_945 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_945 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_946 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_946 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_947 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_947 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_948 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_948 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_949 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_949 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_950 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_950 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_951 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_951 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_952 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_952 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_953 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3b9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_953 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_954 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ba == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_954 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_955 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3bb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_955 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_956 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3bc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_956 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_957 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3bd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_957 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_958 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3be == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_958 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_959 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3bf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_959 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_960 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_960 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_961 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_961 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_962 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_962 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_963 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_963 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_964 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_964 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_965 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_965 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_966 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_966 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_967 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_967 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_968 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_968 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_969 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3c9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_969 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_970 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ca == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_970 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_971 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3cb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_971 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_972 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3cc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_972 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_973 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3cd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_973 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_974 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ce == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_974 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_975 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3cf == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_975 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_976 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_976 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_977 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_977 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_978 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_978 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_979 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_979 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_980 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_980 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_981 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_981 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_982 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_982 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_983 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_983 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_984 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_984 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_985 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3d9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_985 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_986 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3da == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_986 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_987 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3db == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_987 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_988 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3dc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_988 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_989 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3dd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_989 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_990 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3de == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_990 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_991 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3df == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_991 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_992 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_992 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_993 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_993 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_994 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_994 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_995 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_995 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_996 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_996 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_997 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_997 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_998 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_998 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_999 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_999 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1000 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1000 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1001 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3e9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1001 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1002 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ea == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1002 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1003 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3eb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1003 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1004 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ec == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1004 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1005 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ed == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1005 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1006 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ee == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1006 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1007 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ef == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1007 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1008 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f0 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1008 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1009 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f1 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1009 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1010 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f2 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1010 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1011 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f3 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1011 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1012 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f4 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1012 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1013 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f5 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1013 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1014 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f6 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1014 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1015 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f7 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1015 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1016 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f8 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1016 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1017 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3f9 == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1017 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1018 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3fa == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1018 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1019 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3fb == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1019 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1020 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3fc == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1020 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1021 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3fd == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1021 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1022 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3fe == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1022 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
    if (reset) begin // @[OuterBuffer.scala 20:24]
      buffer_1023 <= 16'h0; // @[OuterBuffer.scala 20:24]
    end else if (io_BankIO_Enable) begin // @[OuterBuffer.scala 23:37]
      if (~io_BankIO_ReadWrite) begin // @[OuterBuffer.scala 24:43]
        if (10'h3ff == io_BankIO_DataAddr) begin // @[OuterBuffer.scala 25:34]
          buffer_1023 <= io_BankIO_DataIn; // @[OuterBuffer.scala 25:34]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buffer_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  buffer_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  buffer_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  buffer_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  buffer_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  buffer_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  buffer_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  buffer_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  buffer_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_32 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_33 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  buffer_34 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  buffer_35 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  buffer_36 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_37 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_38 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  buffer_39 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_40 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  buffer_41 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  buffer_42 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_43 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  buffer_44 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_45 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_46 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  buffer_47 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  buffer_48 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  buffer_49 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  buffer_50 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  buffer_51 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  buffer_52 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  buffer_53 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  buffer_54 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  buffer_55 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  buffer_56 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  buffer_57 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  buffer_58 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  buffer_59 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  buffer_60 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  buffer_61 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  buffer_62 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  buffer_63 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  buffer_64 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  buffer_65 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  buffer_66 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  buffer_67 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  buffer_68 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  buffer_69 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  buffer_70 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  buffer_71 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  buffer_72 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  buffer_73 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  buffer_74 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  buffer_75 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  buffer_76 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  buffer_77 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  buffer_78 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  buffer_79 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  buffer_80 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  buffer_81 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  buffer_82 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  buffer_83 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  buffer_84 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  buffer_85 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  buffer_86 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  buffer_87 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  buffer_88 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  buffer_89 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  buffer_90 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  buffer_91 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  buffer_92 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  buffer_93 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  buffer_94 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  buffer_95 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  buffer_96 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  buffer_97 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  buffer_98 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  buffer_99 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  buffer_100 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  buffer_101 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  buffer_102 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  buffer_103 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  buffer_104 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  buffer_105 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  buffer_106 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  buffer_107 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  buffer_108 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  buffer_109 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  buffer_110 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  buffer_111 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  buffer_112 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  buffer_113 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  buffer_114 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  buffer_115 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  buffer_116 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  buffer_117 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  buffer_118 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  buffer_119 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  buffer_120 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  buffer_121 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  buffer_122 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  buffer_123 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  buffer_124 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  buffer_125 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  buffer_126 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  buffer_127 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  buffer_128 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  buffer_129 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  buffer_130 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  buffer_131 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  buffer_132 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  buffer_133 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  buffer_134 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  buffer_135 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  buffer_136 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  buffer_137 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  buffer_138 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  buffer_139 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  buffer_140 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  buffer_141 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  buffer_142 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  buffer_143 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  buffer_144 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  buffer_145 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  buffer_146 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  buffer_147 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  buffer_148 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  buffer_149 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  buffer_150 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  buffer_151 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  buffer_152 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  buffer_153 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  buffer_154 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  buffer_155 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  buffer_156 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  buffer_157 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  buffer_158 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  buffer_159 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  buffer_160 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  buffer_161 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  buffer_162 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  buffer_163 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  buffer_164 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  buffer_165 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  buffer_166 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  buffer_167 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  buffer_168 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  buffer_169 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  buffer_170 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  buffer_171 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  buffer_172 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  buffer_173 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  buffer_174 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  buffer_175 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  buffer_176 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  buffer_177 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  buffer_178 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  buffer_179 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  buffer_180 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  buffer_181 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  buffer_182 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  buffer_183 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  buffer_184 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  buffer_185 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  buffer_186 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  buffer_187 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  buffer_188 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  buffer_189 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  buffer_190 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  buffer_191 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  buffer_192 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  buffer_193 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  buffer_194 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  buffer_195 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  buffer_196 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  buffer_197 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  buffer_198 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  buffer_199 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  buffer_200 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  buffer_201 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  buffer_202 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  buffer_203 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  buffer_204 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  buffer_205 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  buffer_206 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  buffer_207 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  buffer_208 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  buffer_209 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  buffer_210 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  buffer_211 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  buffer_212 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  buffer_213 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  buffer_214 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  buffer_215 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  buffer_216 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  buffer_217 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  buffer_218 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  buffer_219 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  buffer_220 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  buffer_221 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  buffer_222 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  buffer_223 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  buffer_224 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  buffer_225 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  buffer_226 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  buffer_227 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  buffer_228 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  buffer_229 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  buffer_230 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  buffer_231 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  buffer_232 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  buffer_233 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  buffer_234 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  buffer_235 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  buffer_236 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  buffer_237 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  buffer_238 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  buffer_239 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  buffer_240 = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  buffer_241 = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  buffer_242 = _RAND_242[15:0];
  _RAND_243 = {1{`RANDOM}};
  buffer_243 = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  buffer_244 = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  buffer_245 = _RAND_245[15:0];
  _RAND_246 = {1{`RANDOM}};
  buffer_246 = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  buffer_247 = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  buffer_248 = _RAND_248[15:0];
  _RAND_249 = {1{`RANDOM}};
  buffer_249 = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  buffer_250 = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  buffer_251 = _RAND_251[15:0];
  _RAND_252 = {1{`RANDOM}};
  buffer_252 = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  buffer_253 = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  buffer_254 = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  buffer_255 = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  buffer_256 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  buffer_257 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  buffer_258 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  buffer_259 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  buffer_260 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  buffer_261 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  buffer_262 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  buffer_263 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  buffer_264 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  buffer_265 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  buffer_266 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  buffer_267 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  buffer_268 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  buffer_269 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  buffer_270 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  buffer_271 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  buffer_272 = _RAND_272[15:0];
  _RAND_273 = {1{`RANDOM}};
  buffer_273 = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  buffer_274 = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  buffer_275 = _RAND_275[15:0];
  _RAND_276 = {1{`RANDOM}};
  buffer_276 = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  buffer_277 = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  buffer_278 = _RAND_278[15:0];
  _RAND_279 = {1{`RANDOM}};
  buffer_279 = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  buffer_280 = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  buffer_281 = _RAND_281[15:0];
  _RAND_282 = {1{`RANDOM}};
  buffer_282 = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  buffer_283 = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  buffer_284 = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  buffer_285 = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  buffer_286 = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  buffer_287 = _RAND_287[15:0];
  _RAND_288 = {1{`RANDOM}};
  buffer_288 = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  buffer_289 = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  buffer_290 = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  buffer_291 = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  buffer_292 = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  buffer_293 = _RAND_293[15:0];
  _RAND_294 = {1{`RANDOM}};
  buffer_294 = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  buffer_295 = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  buffer_296 = _RAND_296[15:0];
  _RAND_297 = {1{`RANDOM}};
  buffer_297 = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  buffer_298 = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  buffer_299 = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  buffer_300 = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  buffer_301 = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  buffer_302 = _RAND_302[15:0];
  _RAND_303 = {1{`RANDOM}};
  buffer_303 = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  buffer_304 = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  buffer_305 = _RAND_305[15:0];
  _RAND_306 = {1{`RANDOM}};
  buffer_306 = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  buffer_307 = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  buffer_308 = _RAND_308[15:0];
  _RAND_309 = {1{`RANDOM}};
  buffer_309 = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  buffer_310 = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  buffer_311 = _RAND_311[15:0];
  _RAND_312 = {1{`RANDOM}};
  buffer_312 = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  buffer_313 = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  buffer_314 = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  buffer_315 = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  buffer_316 = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  buffer_317 = _RAND_317[15:0];
  _RAND_318 = {1{`RANDOM}};
  buffer_318 = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  buffer_319 = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  buffer_320 = _RAND_320[15:0];
  _RAND_321 = {1{`RANDOM}};
  buffer_321 = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  buffer_322 = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  buffer_323 = _RAND_323[15:0];
  _RAND_324 = {1{`RANDOM}};
  buffer_324 = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  buffer_325 = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  buffer_326 = _RAND_326[15:0];
  _RAND_327 = {1{`RANDOM}};
  buffer_327 = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  buffer_328 = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  buffer_329 = _RAND_329[15:0];
  _RAND_330 = {1{`RANDOM}};
  buffer_330 = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  buffer_331 = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  buffer_332 = _RAND_332[15:0];
  _RAND_333 = {1{`RANDOM}};
  buffer_333 = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  buffer_334 = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  buffer_335 = _RAND_335[15:0];
  _RAND_336 = {1{`RANDOM}};
  buffer_336 = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  buffer_337 = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  buffer_338 = _RAND_338[15:0];
  _RAND_339 = {1{`RANDOM}};
  buffer_339 = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  buffer_340 = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  buffer_341 = _RAND_341[15:0];
  _RAND_342 = {1{`RANDOM}};
  buffer_342 = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  buffer_343 = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  buffer_344 = _RAND_344[15:0];
  _RAND_345 = {1{`RANDOM}};
  buffer_345 = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  buffer_346 = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  buffer_347 = _RAND_347[15:0];
  _RAND_348 = {1{`RANDOM}};
  buffer_348 = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  buffer_349 = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  buffer_350 = _RAND_350[15:0];
  _RAND_351 = {1{`RANDOM}};
  buffer_351 = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  buffer_352 = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  buffer_353 = _RAND_353[15:0];
  _RAND_354 = {1{`RANDOM}};
  buffer_354 = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  buffer_355 = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  buffer_356 = _RAND_356[15:0];
  _RAND_357 = {1{`RANDOM}};
  buffer_357 = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  buffer_358 = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  buffer_359 = _RAND_359[15:0];
  _RAND_360 = {1{`RANDOM}};
  buffer_360 = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  buffer_361 = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  buffer_362 = _RAND_362[15:0];
  _RAND_363 = {1{`RANDOM}};
  buffer_363 = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  buffer_364 = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  buffer_365 = _RAND_365[15:0];
  _RAND_366 = {1{`RANDOM}};
  buffer_366 = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  buffer_367 = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  buffer_368 = _RAND_368[15:0];
  _RAND_369 = {1{`RANDOM}};
  buffer_369 = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  buffer_370 = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  buffer_371 = _RAND_371[15:0];
  _RAND_372 = {1{`RANDOM}};
  buffer_372 = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  buffer_373 = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  buffer_374 = _RAND_374[15:0];
  _RAND_375 = {1{`RANDOM}};
  buffer_375 = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  buffer_376 = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  buffer_377 = _RAND_377[15:0];
  _RAND_378 = {1{`RANDOM}};
  buffer_378 = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  buffer_379 = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  buffer_380 = _RAND_380[15:0];
  _RAND_381 = {1{`RANDOM}};
  buffer_381 = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  buffer_382 = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  buffer_383 = _RAND_383[15:0];
  _RAND_384 = {1{`RANDOM}};
  buffer_384 = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  buffer_385 = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  buffer_386 = _RAND_386[15:0];
  _RAND_387 = {1{`RANDOM}};
  buffer_387 = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  buffer_388 = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  buffer_389 = _RAND_389[15:0];
  _RAND_390 = {1{`RANDOM}};
  buffer_390 = _RAND_390[15:0];
  _RAND_391 = {1{`RANDOM}};
  buffer_391 = _RAND_391[15:0];
  _RAND_392 = {1{`RANDOM}};
  buffer_392 = _RAND_392[15:0];
  _RAND_393 = {1{`RANDOM}};
  buffer_393 = _RAND_393[15:0];
  _RAND_394 = {1{`RANDOM}};
  buffer_394 = _RAND_394[15:0];
  _RAND_395 = {1{`RANDOM}};
  buffer_395 = _RAND_395[15:0];
  _RAND_396 = {1{`RANDOM}};
  buffer_396 = _RAND_396[15:0];
  _RAND_397 = {1{`RANDOM}};
  buffer_397 = _RAND_397[15:0];
  _RAND_398 = {1{`RANDOM}};
  buffer_398 = _RAND_398[15:0];
  _RAND_399 = {1{`RANDOM}};
  buffer_399 = _RAND_399[15:0];
  _RAND_400 = {1{`RANDOM}};
  buffer_400 = _RAND_400[15:0];
  _RAND_401 = {1{`RANDOM}};
  buffer_401 = _RAND_401[15:0];
  _RAND_402 = {1{`RANDOM}};
  buffer_402 = _RAND_402[15:0];
  _RAND_403 = {1{`RANDOM}};
  buffer_403 = _RAND_403[15:0];
  _RAND_404 = {1{`RANDOM}};
  buffer_404 = _RAND_404[15:0];
  _RAND_405 = {1{`RANDOM}};
  buffer_405 = _RAND_405[15:0];
  _RAND_406 = {1{`RANDOM}};
  buffer_406 = _RAND_406[15:0];
  _RAND_407 = {1{`RANDOM}};
  buffer_407 = _RAND_407[15:0];
  _RAND_408 = {1{`RANDOM}};
  buffer_408 = _RAND_408[15:0];
  _RAND_409 = {1{`RANDOM}};
  buffer_409 = _RAND_409[15:0];
  _RAND_410 = {1{`RANDOM}};
  buffer_410 = _RAND_410[15:0];
  _RAND_411 = {1{`RANDOM}};
  buffer_411 = _RAND_411[15:0];
  _RAND_412 = {1{`RANDOM}};
  buffer_412 = _RAND_412[15:0];
  _RAND_413 = {1{`RANDOM}};
  buffer_413 = _RAND_413[15:0];
  _RAND_414 = {1{`RANDOM}};
  buffer_414 = _RAND_414[15:0];
  _RAND_415 = {1{`RANDOM}};
  buffer_415 = _RAND_415[15:0];
  _RAND_416 = {1{`RANDOM}};
  buffer_416 = _RAND_416[15:0];
  _RAND_417 = {1{`RANDOM}};
  buffer_417 = _RAND_417[15:0];
  _RAND_418 = {1{`RANDOM}};
  buffer_418 = _RAND_418[15:0];
  _RAND_419 = {1{`RANDOM}};
  buffer_419 = _RAND_419[15:0];
  _RAND_420 = {1{`RANDOM}};
  buffer_420 = _RAND_420[15:0];
  _RAND_421 = {1{`RANDOM}};
  buffer_421 = _RAND_421[15:0];
  _RAND_422 = {1{`RANDOM}};
  buffer_422 = _RAND_422[15:0];
  _RAND_423 = {1{`RANDOM}};
  buffer_423 = _RAND_423[15:0];
  _RAND_424 = {1{`RANDOM}};
  buffer_424 = _RAND_424[15:0];
  _RAND_425 = {1{`RANDOM}};
  buffer_425 = _RAND_425[15:0];
  _RAND_426 = {1{`RANDOM}};
  buffer_426 = _RAND_426[15:0];
  _RAND_427 = {1{`RANDOM}};
  buffer_427 = _RAND_427[15:0];
  _RAND_428 = {1{`RANDOM}};
  buffer_428 = _RAND_428[15:0];
  _RAND_429 = {1{`RANDOM}};
  buffer_429 = _RAND_429[15:0];
  _RAND_430 = {1{`RANDOM}};
  buffer_430 = _RAND_430[15:0];
  _RAND_431 = {1{`RANDOM}};
  buffer_431 = _RAND_431[15:0];
  _RAND_432 = {1{`RANDOM}};
  buffer_432 = _RAND_432[15:0];
  _RAND_433 = {1{`RANDOM}};
  buffer_433 = _RAND_433[15:0];
  _RAND_434 = {1{`RANDOM}};
  buffer_434 = _RAND_434[15:0];
  _RAND_435 = {1{`RANDOM}};
  buffer_435 = _RAND_435[15:0];
  _RAND_436 = {1{`RANDOM}};
  buffer_436 = _RAND_436[15:0];
  _RAND_437 = {1{`RANDOM}};
  buffer_437 = _RAND_437[15:0];
  _RAND_438 = {1{`RANDOM}};
  buffer_438 = _RAND_438[15:0];
  _RAND_439 = {1{`RANDOM}};
  buffer_439 = _RAND_439[15:0];
  _RAND_440 = {1{`RANDOM}};
  buffer_440 = _RAND_440[15:0];
  _RAND_441 = {1{`RANDOM}};
  buffer_441 = _RAND_441[15:0];
  _RAND_442 = {1{`RANDOM}};
  buffer_442 = _RAND_442[15:0];
  _RAND_443 = {1{`RANDOM}};
  buffer_443 = _RAND_443[15:0];
  _RAND_444 = {1{`RANDOM}};
  buffer_444 = _RAND_444[15:0];
  _RAND_445 = {1{`RANDOM}};
  buffer_445 = _RAND_445[15:0];
  _RAND_446 = {1{`RANDOM}};
  buffer_446 = _RAND_446[15:0];
  _RAND_447 = {1{`RANDOM}};
  buffer_447 = _RAND_447[15:0];
  _RAND_448 = {1{`RANDOM}};
  buffer_448 = _RAND_448[15:0];
  _RAND_449 = {1{`RANDOM}};
  buffer_449 = _RAND_449[15:0];
  _RAND_450 = {1{`RANDOM}};
  buffer_450 = _RAND_450[15:0];
  _RAND_451 = {1{`RANDOM}};
  buffer_451 = _RAND_451[15:0];
  _RAND_452 = {1{`RANDOM}};
  buffer_452 = _RAND_452[15:0];
  _RAND_453 = {1{`RANDOM}};
  buffer_453 = _RAND_453[15:0];
  _RAND_454 = {1{`RANDOM}};
  buffer_454 = _RAND_454[15:0];
  _RAND_455 = {1{`RANDOM}};
  buffer_455 = _RAND_455[15:0];
  _RAND_456 = {1{`RANDOM}};
  buffer_456 = _RAND_456[15:0];
  _RAND_457 = {1{`RANDOM}};
  buffer_457 = _RAND_457[15:0];
  _RAND_458 = {1{`RANDOM}};
  buffer_458 = _RAND_458[15:0];
  _RAND_459 = {1{`RANDOM}};
  buffer_459 = _RAND_459[15:0];
  _RAND_460 = {1{`RANDOM}};
  buffer_460 = _RAND_460[15:0];
  _RAND_461 = {1{`RANDOM}};
  buffer_461 = _RAND_461[15:0];
  _RAND_462 = {1{`RANDOM}};
  buffer_462 = _RAND_462[15:0];
  _RAND_463 = {1{`RANDOM}};
  buffer_463 = _RAND_463[15:0];
  _RAND_464 = {1{`RANDOM}};
  buffer_464 = _RAND_464[15:0];
  _RAND_465 = {1{`RANDOM}};
  buffer_465 = _RAND_465[15:0];
  _RAND_466 = {1{`RANDOM}};
  buffer_466 = _RAND_466[15:0];
  _RAND_467 = {1{`RANDOM}};
  buffer_467 = _RAND_467[15:0];
  _RAND_468 = {1{`RANDOM}};
  buffer_468 = _RAND_468[15:0];
  _RAND_469 = {1{`RANDOM}};
  buffer_469 = _RAND_469[15:0];
  _RAND_470 = {1{`RANDOM}};
  buffer_470 = _RAND_470[15:0];
  _RAND_471 = {1{`RANDOM}};
  buffer_471 = _RAND_471[15:0];
  _RAND_472 = {1{`RANDOM}};
  buffer_472 = _RAND_472[15:0];
  _RAND_473 = {1{`RANDOM}};
  buffer_473 = _RAND_473[15:0];
  _RAND_474 = {1{`RANDOM}};
  buffer_474 = _RAND_474[15:0];
  _RAND_475 = {1{`RANDOM}};
  buffer_475 = _RAND_475[15:0];
  _RAND_476 = {1{`RANDOM}};
  buffer_476 = _RAND_476[15:0];
  _RAND_477 = {1{`RANDOM}};
  buffer_477 = _RAND_477[15:0];
  _RAND_478 = {1{`RANDOM}};
  buffer_478 = _RAND_478[15:0];
  _RAND_479 = {1{`RANDOM}};
  buffer_479 = _RAND_479[15:0];
  _RAND_480 = {1{`RANDOM}};
  buffer_480 = _RAND_480[15:0];
  _RAND_481 = {1{`RANDOM}};
  buffer_481 = _RAND_481[15:0];
  _RAND_482 = {1{`RANDOM}};
  buffer_482 = _RAND_482[15:0];
  _RAND_483 = {1{`RANDOM}};
  buffer_483 = _RAND_483[15:0];
  _RAND_484 = {1{`RANDOM}};
  buffer_484 = _RAND_484[15:0];
  _RAND_485 = {1{`RANDOM}};
  buffer_485 = _RAND_485[15:0];
  _RAND_486 = {1{`RANDOM}};
  buffer_486 = _RAND_486[15:0];
  _RAND_487 = {1{`RANDOM}};
  buffer_487 = _RAND_487[15:0];
  _RAND_488 = {1{`RANDOM}};
  buffer_488 = _RAND_488[15:0];
  _RAND_489 = {1{`RANDOM}};
  buffer_489 = _RAND_489[15:0];
  _RAND_490 = {1{`RANDOM}};
  buffer_490 = _RAND_490[15:0];
  _RAND_491 = {1{`RANDOM}};
  buffer_491 = _RAND_491[15:0];
  _RAND_492 = {1{`RANDOM}};
  buffer_492 = _RAND_492[15:0];
  _RAND_493 = {1{`RANDOM}};
  buffer_493 = _RAND_493[15:0];
  _RAND_494 = {1{`RANDOM}};
  buffer_494 = _RAND_494[15:0];
  _RAND_495 = {1{`RANDOM}};
  buffer_495 = _RAND_495[15:0];
  _RAND_496 = {1{`RANDOM}};
  buffer_496 = _RAND_496[15:0];
  _RAND_497 = {1{`RANDOM}};
  buffer_497 = _RAND_497[15:0];
  _RAND_498 = {1{`RANDOM}};
  buffer_498 = _RAND_498[15:0];
  _RAND_499 = {1{`RANDOM}};
  buffer_499 = _RAND_499[15:0];
  _RAND_500 = {1{`RANDOM}};
  buffer_500 = _RAND_500[15:0];
  _RAND_501 = {1{`RANDOM}};
  buffer_501 = _RAND_501[15:0];
  _RAND_502 = {1{`RANDOM}};
  buffer_502 = _RAND_502[15:0];
  _RAND_503 = {1{`RANDOM}};
  buffer_503 = _RAND_503[15:0];
  _RAND_504 = {1{`RANDOM}};
  buffer_504 = _RAND_504[15:0];
  _RAND_505 = {1{`RANDOM}};
  buffer_505 = _RAND_505[15:0];
  _RAND_506 = {1{`RANDOM}};
  buffer_506 = _RAND_506[15:0];
  _RAND_507 = {1{`RANDOM}};
  buffer_507 = _RAND_507[15:0];
  _RAND_508 = {1{`RANDOM}};
  buffer_508 = _RAND_508[15:0];
  _RAND_509 = {1{`RANDOM}};
  buffer_509 = _RAND_509[15:0];
  _RAND_510 = {1{`RANDOM}};
  buffer_510 = _RAND_510[15:0];
  _RAND_511 = {1{`RANDOM}};
  buffer_511 = _RAND_511[15:0];
  _RAND_512 = {1{`RANDOM}};
  buffer_512 = _RAND_512[15:0];
  _RAND_513 = {1{`RANDOM}};
  buffer_513 = _RAND_513[15:0];
  _RAND_514 = {1{`RANDOM}};
  buffer_514 = _RAND_514[15:0];
  _RAND_515 = {1{`RANDOM}};
  buffer_515 = _RAND_515[15:0];
  _RAND_516 = {1{`RANDOM}};
  buffer_516 = _RAND_516[15:0];
  _RAND_517 = {1{`RANDOM}};
  buffer_517 = _RAND_517[15:0];
  _RAND_518 = {1{`RANDOM}};
  buffer_518 = _RAND_518[15:0];
  _RAND_519 = {1{`RANDOM}};
  buffer_519 = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  buffer_520 = _RAND_520[15:0];
  _RAND_521 = {1{`RANDOM}};
  buffer_521 = _RAND_521[15:0];
  _RAND_522 = {1{`RANDOM}};
  buffer_522 = _RAND_522[15:0];
  _RAND_523 = {1{`RANDOM}};
  buffer_523 = _RAND_523[15:0];
  _RAND_524 = {1{`RANDOM}};
  buffer_524 = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  buffer_525 = _RAND_525[15:0];
  _RAND_526 = {1{`RANDOM}};
  buffer_526 = _RAND_526[15:0];
  _RAND_527 = {1{`RANDOM}};
  buffer_527 = _RAND_527[15:0];
  _RAND_528 = {1{`RANDOM}};
  buffer_528 = _RAND_528[15:0];
  _RAND_529 = {1{`RANDOM}};
  buffer_529 = _RAND_529[15:0];
  _RAND_530 = {1{`RANDOM}};
  buffer_530 = _RAND_530[15:0];
  _RAND_531 = {1{`RANDOM}};
  buffer_531 = _RAND_531[15:0];
  _RAND_532 = {1{`RANDOM}};
  buffer_532 = _RAND_532[15:0];
  _RAND_533 = {1{`RANDOM}};
  buffer_533 = _RAND_533[15:0];
  _RAND_534 = {1{`RANDOM}};
  buffer_534 = _RAND_534[15:0];
  _RAND_535 = {1{`RANDOM}};
  buffer_535 = _RAND_535[15:0];
  _RAND_536 = {1{`RANDOM}};
  buffer_536 = _RAND_536[15:0];
  _RAND_537 = {1{`RANDOM}};
  buffer_537 = _RAND_537[15:0];
  _RAND_538 = {1{`RANDOM}};
  buffer_538 = _RAND_538[15:0];
  _RAND_539 = {1{`RANDOM}};
  buffer_539 = _RAND_539[15:0];
  _RAND_540 = {1{`RANDOM}};
  buffer_540 = _RAND_540[15:0];
  _RAND_541 = {1{`RANDOM}};
  buffer_541 = _RAND_541[15:0];
  _RAND_542 = {1{`RANDOM}};
  buffer_542 = _RAND_542[15:0];
  _RAND_543 = {1{`RANDOM}};
  buffer_543 = _RAND_543[15:0];
  _RAND_544 = {1{`RANDOM}};
  buffer_544 = _RAND_544[15:0];
  _RAND_545 = {1{`RANDOM}};
  buffer_545 = _RAND_545[15:0];
  _RAND_546 = {1{`RANDOM}};
  buffer_546 = _RAND_546[15:0];
  _RAND_547 = {1{`RANDOM}};
  buffer_547 = _RAND_547[15:0];
  _RAND_548 = {1{`RANDOM}};
  buffer_548 = _RAND_548[15:0];
  _RAND_549 = {1{`RANDOM}};
  buffer_549 = _RAND_549[15:0];
  _RAND_550 = {1{`RANDOM}};
  buffer_550 = _RAND_550[15:0];
  _RAND_551 = {1{`RANDOM}};
  buffer_551 = _RAND_551[15:0];
  _RAND_552 = {1{`RANDOM}};
  buffer_552 = _RAND_552[15:0];
  _RAND_553 = {1{`RANDOM}};
  buffer_553 = _RAND_553[15:0];
  _RAND_554 = {1{`RANDOM}};
  buffer_554 = _RAND_554[15:0];
  _RAND_555 = {1{`RANDOM}};
  buffer_555 = _RAND_555[15:0];
  _RAND_556 = {1{`RANDOM}};
  buffer_556 = _RAND_556[15:0];
  _RAND_557 = {1{`RANDOM}};
  buffer_557 = _RAND_557[15:0];
  _RAND_558 = {1{`RANDOM}};
  buffer_558 = _RAND_558[15:0];
  _RAND_559 = {1{`RANDOM}};
  buffer_559 = _RAND_559[15:0];
  _RAND_560 = {1{`RANDOM}};
  buffer_560 = _RAND_560[15:0];
  _RAND_561 = {1{`RANDOM}};
  buffer_561 = _RAND_561[15:0];
  _RAND_562 = {1{`RANDOM}};
  buffer_562 = _RAND_562[15:0];
  _RAND_563 = {1{`RANDOM}};
  buffer_563 = _RAND_563[15:0];
  _RAND_564 = {1{`RANDOM}};
  buffer_564 = _RAND_564[15:0];
  _RAND_565 = {1{`RANDOM}};
  buffer_565 = _RAND_565[15:0];
  _RAND_566 = {1{`RANDOM}};
  buffer_566 = _RAND_566[15:0];
  _RAND_567 = {1{`RANDOM}};
  buffer_567 = _RAND_567[15:0];
  _RAND_568 = {1{`RANDOM}};
  buffer_568 = _RAND_568[15:0];
  _RAND_569 = {1{`RANDOM}};
  buffer_569 = _RAND_569[15:0];
  _RAND_570 = {1{`RANDOM}};
  buffer_570 = _RAND_570[15:0];
  _RAND_571 = {1{`RANDOM}};
  buffer_571 = _RAND_571[15:0];
  _RAND_572 = {1{`RANDOM}};
  buffer_572 = _RAND_572[15:0];
  _RAND_573 = {1{`RANDOM}};
  buffer_573 = _RAND_573[15:0];
  _RAND_574 = {1{`RANDOM}};
  buffer_574 = _RAND_574[15:0];
  _RAND_575 = {1{`RANDOM}};
  buffer_575 = _RAND_575[15:0];
  _RAND_576 = {1{`RANDOM}};
  buffer_576 = _RAND_576[15:0];
  _RAND_577 = {1{`RANDOM}};
  buffer_577 = _RAND_577[15:0];
  _RAND_578 = {1{`RANDOM}};
  buffer_578 = _RAND_578[15:0];
  _RAND_579 = {1{`RANDOM}};
  buffer_579 = _RAND_579[15:0];
  _RAND_580 = {1{`RANDOM}};
  buffer_580 = _RAND_580[15:0];
  _RAND_581 = {1{`RANDOM}};
  buffer_581 = _RAND_581[15:0];
  _RAND_582 = {1{`RANDOM}};
  buffer_582 = _RAND_582[15:0];
  _RAND_583 = {1{`RANDOM}};
  buffer_583 = _RAND_583[15:0];
  _RAND_584 = {1{`RANDOM}};
  buffer_584 = _RAND_584[15:0];
  _RAND_585 = {1{`RANDOM}};
  buffer_585 = _RAND_585[15:0];
  _RAND_586 = {1{`RANDOM}};
  buffer_586 = _RAND_586[15:0];
  _RAND_587 = {1{`RANDOM}};
  buffer_587 = _RAND_587[15:0];
  _RAND_588 = {1{`RANDOM}};
  buffer_588 = _RAND_588[15:0];
  _RAND_589 = {1{`RANDOM}};
  buffer_589 = _RAND_589[15:0];
  _RAND_590 = {1{`RANDOM}};
  buffer_590 = _RAND_590[15:0];
  _RAND_591 = {1{`RANDOM}};
  buffer_591 = _RAND_591[15:0];
  _RAND_592 = {1{`RANDOM}};
  buffer_592 = _RAND_592[15:0];
  _RAND_593 = {1{`RANDOM}};
  buffer_593 = _RAND_593[15:0];
  _RAND_594 = {1{`RANDOM}};
  buffer_594 = _RAND_594[15:0];
  _RAND_595 = {1{`RANDOM}};
  buffer_595 = _RAND_595[15:0];
  _RAND_596 = {1{`RANDOM}};
  buffer_596 = _RAND_596[15:0];
  _RAND_597 = {1{`RANDOM}};
  buffer_597 = _RAND_597[15:0];
  _RAND_598 = {1{`RANDOM}};
  buffer_598 = _RAND_598[15:0];
  _RAND_599 = {1{`RANDOM}};
  buffer_599 = _RAND_599[15:0];
  _RAND_600 = {1{`RANDOM}};
  buffer_600 = _RAND_600[15:0];
  _RAND_601 = {1{`RANDOM}};
  buffer_601 = _RAND_601[15:0];
  _RAND_602 = {1{`RANDOM}};
  buffer_602 = _RAND_602[15:0];
  _RAND_603 = {1{`RANDOM}};
  buffer_603 = _RAND_603[15:0];
  _RAND_604 = {1{`RANDOM}};
  buffer_604 = _RAND_604[15:0];
  _RAND_605 = {1{`RANDOM}};
  buffer_605 = _RAND_605[15:0];
  _RAND_606 = {1{`RANDOM}};
  buffer_606 = _RAND_606[15:0];
  _RAND_607 = {1{`RANDOM}};
  buffer_607 = _RAND_607[15:0];
  _RAND_608 = {1{`RANDOM}};
  buffer_608 = _RAND_608[15:0];
  _RAND_609 = {1{`RANDOM}};
  buffer_609 = _RAND_609[15:0];
  _RAND_610 = {1{`RANDOM}};
  buffer_610 = _RAND_610[15:0];
  _RAND_611 = {1{`RANDOM}};
  buffer_611 = _RAND_611[15:0];
  _RAND_612 = {1{`RANDOM}};
  buffer_612 = _RAND_612[15:0];
  _RAND_613 = {1{`RANDOM}};
  buffer_613 = _RAND_613[15:0];
  _RAND_614 = {1{`RANDOM}};
  buffer_614 = _RAND_614[15:0];
  _RAND_615 = {1{`RANDOM}};
  buffer_615 = _RAND_615[15:0];
  _RAND_616 = {1{`RANDOM}};
  buffer_616 = _RAND_616[15:0];
  _RAND_617 = {1{`RANDOM}};
  buffer_617 = _RAND_617[15:0];
  _RAND_618 = {1{`RANDOM}};
  buffer_618 = _RAND_618[15:0];
  _RAND_619 = {1{`RANDOM}};
  buffer_619 = _RAND_619[15:0];
  _RAND_620 = {1{`RANDOM}};
  buffer_620 = _RAND_620[15:0];
  _RAND_621 = {1{`RANDOM}};
  buffer_621 = _RAND_621[15:0];
  _RAND_622 = {1{`RANDOM}};
  buffer_622 = _RAND_622[15:0];
  _RAND_623 = {1{`RANDOM}};
  buffer_623 = _RAND_623[15:0];
  _RAND_624 = {1{`RANDOM}};
  buffer_624 = _RAND_624[15:0];
  _RAND_625 = {1{`RANDOM}};
  buffer_625 = _RAND_625[15:0];
  _RAND_626 = {1{`RANDOM}};
  buffer_626 = _RAND_626[15:0];
  _RAND_627 = {1{`RANDOM}};
  buffer_627 = _RAND_627[15:0];
  _RAND_628 = {1{`RANDOM}};
  buffer_628 = _RAND_628[15:0];
  _RAND_629 = {1{`RANDOM}};
  buffer_629 = _RAND_629[15:0];
  _RAND_630 = {1{`RANDOM}};
  buffer_630 = _RAND_630[15:0];
  _RAND_631 = {1{`RANDOM}};
  buffer_631 = _RAND_631[15:0];
  _RAND_632 = {1{`RANDOM}};
  buffer_632 = _RAND_632[15:0];
  _RAND_633 = {1{`RANDOM}};
  buffer_633 = _RAND_633[15:0];
  _RAND_634 = {1{`RANDOM}};
  buffer_634 = _RAND_634[15:0];
  _RAND_635 = {1{`RANDOM}};
  buffer_635 = _RAND_635[15:0];
  _RAND_636 = {1{`RANDOM}};
  buffer_636 = _RAND_636[15:0];
  _RAND_637 = {1{`RANDOM}};
  buffer_637 = _RAND_637[15:0];
  _RAND_638 = {1{`RANDOM}};
  buffer_638 = _RAND_638[15:0];
  _RAND_639 = {1{`RANDOM}};
  buffer_639 = _RAND_639[15:0];
  _RAND_640 = {1{`RANDOM}};
  buffer_640 = _RAND_640[15:0];
  _RAND_641 = {1{`RANDOM}};
  buffer_641 = _RAND_641[15:0];
  _RAND_642 = {1{`RANDOM}};
  buffer_642 = _RAND_642[15:0];
  _RAND_643 = {1{`RANDOM}};
  buffer_643 = _RAND_643[15:0];
  _RAND_644 = {1{`RANDOM}};
  buffer_644 = _RAND_644[15:0];
  _RAND_645 = {1{`RANDOM}};
  buffer_645 = _RAND_645[15:0];
  _RAND_646 = {1{`RANDOM}};
  buffer_646 = _RAND_646[15:0];
  _RAND_647 = {1{`RANDOM}};
  buffer_647 = _RAND_647[15:0];
  _RAND_648 = {1{`RANDOM}};
  buffer_648 = _RAND_648[15:0];
  _RAND_649 = {1{`RANDOM}};
  buffer_649 = _RAND_649[15:0];
  _RAND_650 = {1{`RANDOM}};
  buffer_650 = _RAND_650[15:0];
  _RAND_651 = {1{`RANDOM}};
  buffer_651 = _RAND_651[15:0];
  _RAND_652 = {1{`RANDOM}};
  buffer_652 = _RAND_652[15:0];
  _RAND_653 = {1{`RANDOM}};
  buffer_653 = _RAND_653[15:0];
  _RAND_654 = {1{`RANDOM}};
  buffer_654 = _RAND_654[15:0];
  _RAND_655 = {1{`RANDOM}};
  buffer_655 = _RAND_655[15:0];
  _RAND_656 = {1{`RANDOM}};
  buffer_656 = _RAND_656[15:0];
  _RAND_657 = {1{`RANDOM}};
  buffer_657 = _RAND_657[15:0];
  _RAND_658 = {1{`RANDOM}};
  buffer_658 = _RAND_658[15:0];
  _RAND_659 = {1{`RANDOM}};
  buffer_659 = _RAND_659[15:0];
  _RAND_660 = {1{`RANDOM}};
  buffer_660 = _RAND_660[15:0];
  _RAND_661 = {1{`RANDOM}};
  buffer_661 = _RAND_661[15:0];
  _RAND_662 = {1{`RANDOM}};
  buffer_662 = _RAND_662[15:0];
  _RAND_663 = {1{`RANDOM}};
  buffer_663 = _RAND_663[15:0];
  _RAND_664 = {1{`RANDOM}};
  buffer_664 = _RAND_664[15:0];
  _RAND_665 = {1{`RANDOM}};
  buffer_665 = _RAND_665[15:0];
  _RAND_666 = {1{`RANDOM}};
  buffer_666 = _RAND_666[15:0];
  _RAND_667 = {1{`RANDOM}};
  buffer_667 = _RAND_667[15:0];
  _RAND_668 = {1{`RANDOM}};
  buffer_668 = _RAND_668[15:0];
  _RAND_669 = {1{`RANDOM}};
  buffer_669 = _RAND_669[15:0];
  _RAND_670 = {1{`RANDOM}};
  buffer_670 = _RAND_670[15:0];
  _RAND_671 = {1{`RANDOM}};
  buffer_671 = _RAND_671[15:0];
  _RAND_672 = {1{`RANDOM}};
  buffer_672 = _RAND_672[15:0];
  _RAND_673 = {1{`RANDOM}};
  buffer_673 = _RAND_673[15:0];
  _RAND_674 = {1{`RANDOM}};
  buffer_674 = _RAND_674[15:0];
  _RAND_675 = {1{`RANDOM}};
  buffer_675 = _RAND_675[15:0];
  _RAND_676 = {1{`RANDOM}};
  buffer_676 = _RAND_676[15:0];
  _RAND_677 = {1{`RANDOM}};
  buffer_677 = _RAND_677[15:0];
  _RAND_678 = {1{`RANDOM}};
  buffer_678 = _RAND_678[15:0];
  _RAND_679 = {1{`RANDOM}};
  buffer_679 = _RAND_679[15:0];
  _RAND_680 = {1{`RANDOM}};
  buffer_680 = _RAND_680[15:0];
  _RAND_681 = {1{`RANDOM}};
  buffer_681 = _RAND_681[15:0];
  _RAND_682 = {1{`RANDOM}};
  buffer_682 = _RAND_682[15:0];
  _RAND_683 = {1{`RANDOM}};
  buffer_683 = _RAND_683[15:0];
  _RAND_684 = {1{`RANDOM}};
  buffer_684 = _RAND_684[15:0];
  _RAND_685 = {1{`RANDOM}};
  buffer_685 = _RAND_685[15:0];
  _RAND_686 = {1{`RANDOM}};
  buffer_686 = _RAND_686[15:0];
  _RAND_687 = {1{`RANDOM}};
  buffer_687 = _RAND_687[15:0];
  _RAND_688 = {1{`RANDOM}};
  buffer_688 = _RAND_688[15:0];
  _RAND_689 = {1{`RANDOM}};
  buffer_689 = _RAND_689[15:0];
  _RAND_690 = {1{`RANDOM}};
  buffer_690 = _RAND_690[15:0];
  _RAND_691 = {1{`RANDOM}};
  buffer_691 = _RAND_691[15:0];
  _RAND_692 = {1{`RANDOM}};
  buffer_692 = _RAND_692[15:0];
  _RAND_693 = {1{`RANDOM}};
  buffer_693 = _RAND_693[15:0];
  _RAND_694 = {1{`RANDOM}};
  buffer_694 = _RAND_694[15:0];
  _RAND_695 = {1{`RANDOM}};
  buffer_695 = _RAND_695[15:0];
  _RAND_696 = {1{`RANDOM}};
  buffer_696 = _RAND_696[15:0];
  _RAND_697 = {1{`RANDOM}};
  buffer_697 = _RAND_697[15:0];
  _RAND_698 = {1{`RANDOM}};
  buffer_698 = _RAND_698[15:0];
  _RAND_699 = {1{`RANDOM}};
  buffer_699 = _RAND_699[15:0];
  _RAND_700 = {1{`RANDOM}};
  buffer_700 = _RAND_700[15:0];
  _RAND_701 = {1{`RANDOM}};
  buffer_701 = _RAND_701[15:0];
  _RAND_702 = {1{`RANDOM}};
  buffer_702 = _RAND_702[15:0];
  _RAND_703 = {1{`RANDOM}};
  buffer_703 = _RAND_703[15:0];
  _RAND_704 = {1{`RANDOM}};
  buffer_704 = _RAND_704[15:0];
  _RAND_705 = {1{`RANDOM}};
  buffer_705 = _RAND_705[15:0];
  _RAND_706 = {1{`RANDOM}};
  buffer_706 = _RAND_706[15:0];
  _RAND_707 = {1{`RANDOM}};
  buffer_707 = _RAND_707[15:0];
  _RAND_708 = {1{`RANDOM}};
  buffer_708 = _RAND_708[15:0];
  _RAND_709 = {1{`RANDOM}};
  buffer_709 = _RAND_709[15:0];
  _RAND_710 = {1{`RANDOM}};
  buffer_710 = _RAND_710[15:0];
  _RAND_711 = {1{`RANDOM}};
  buffer_711 = _RAND_711[15:0];
  _RAND_712 = {1{`RANDOM}};
  buffer_712 = _RAND_712[15:0];
  _RAND_713 = {1{`RANDOM}};
  buffer_713 = _RAND_713[15:0];
  _RAND_714 = {1{`RANDOM}};
  buffer_714 = _RAND_714[15:0];
  _RAND_715 = {1{`RANDOM}};
  buffer_715 = _RAND_715[15:0];
  _RAND_716 = {1{`RANDOM}};
  buffer_716 = _RAND_716[15:0];
  _RAND_717 = {1{`RANDOM}};
  buffer_717 = _RAND_717[15:0];
  _RAND_718 = {1{`RANDOM}};
  buffer_718 = _RAND_718[15:0];
  _RAND_719 = {1{`RANDOM}};
  buffer_719 = _RAND_719[15:0];
  _RAND_720 = {1{`RANDOM}};
  buffer_720 = _RAND_720[15:0];
  _RAND_721 = {1{`RANDOM}};
  buffer_721 = _RAND_721[15:0];
  _RAND_722 = {1{`RANDOM}};
  buffer_722 = _RAND_722[15:0];
  _RAND_723 = {1{`RANDOM}};
  buffer_723 = _RAND_723[15:0];
  _RAND_724 = {1{`RANDOM}};
  buffer_724 = _RAND_724[15:0];
  _RAND_725 = {1{`RANDOM}};
  buffer_725 = _RAND_725[15:0];
  _RAND_726 = {1{`RANDOM}};
  buffer_726 = _RAND_726[15:0];
  _RAND_727 = {1{`RANDOM}};
  buffer_727 = _RAND_727[15:0];
  _RAND_728 = {1{`RANDOM}};
  buffer_728 = _RAND_728[15:0];
  _RAND_729 = {1{`RANDOM}};
  buffer_729 = _RAND_729[15:0];
  _RAND_730 = {1{`RANDOM}};
  buffer_730 = _RAND_730[15:0];
  _RAND_731 = {1{`RANDOM}};
  buffer_731 = _RAND_731[15:0];
  _RAND_732 = {1{`RANDOM}};
  buffer_732 = _RAND_732[15:0];
  _RAND_733 = {1{`RANDOM}};
  buffer_733 = _RAND_733[15:0];
  _RAND_734 = {1{`RANDOM}};
  buffer_734 = _RAND_734[15:0];
  _RAND_735 = {1{`RANDOM}};
  buffer_735 = _RAND_735[15:0];
  _RAND_736 = {1{`RANDOM}};
  buffer_736 = _RAND_736[15:0];
  _RAND_737 = {1{`RANDOM}};
  buffer_737 = _RAND_737[15:0];
  _RAND_738 = {1{`RANDOM}};
  buffer_738 = _RAND_738[15:0];
  _RAND_739 = {1{`RANDOM}};
  buffer_739 = _RAND_739[15:0];
  _RAND_740 = {1{`RANDOM}};
  buffer_740 = _RAND_740[15:0];
  _RAND_741 = {1{`RANDOM}};
  buffer_741 = _RAND_741[15:0];
  _RAND_742 = {1{`RANDOM}};
  buffer_742 = _RAND_742[15:0];
  _RAND_743 = {1{`RANDOM}};
  buffer_743 = _RAND_743[15:0];
  _RAND_744 = {1{`RANDOM}};
  buffer_744 = _RAND_744[15:0];
  _RAND_745 = {1{`RANDOM}};
  buffer_745 = _RAND_745[15:0];
  _RAND_746 = {1{`RANDOM}};
  buffer_746 = _RAND_746[15:0];
  _RAND_747 = {1{`RANDOM}};
  buffer_747 = _RAND_747[15:0];
  _RAND_748 = {1{`RANDOM}};
  buffer_748 = _RAND_748[15:0];
  _RAND_749 = {1{`RANDOM}};
  buffer_749 = _RAND_749[15:0];
  _RAND_750 = {1{`RANDOM}};
  buffer_750 = _RAND_750[15:0];
  _RAND_751 = {1{`RANDOM}};
  buffer_751 = _RAND_751[15:0];
  _RAND_752 = {1{`RANDOM}};
  buffer_752 = _RAND_752[15:0];
  _RAND_753 = {1{`RANDOM}};
  buffer_753 = _RAND_753[15:0];
  _RAND_754 = {1{`RANDOM}};
  buffer_754 = _RAND_754[15:0];
  _RAND_755 = {1{`RANDOM}};
  buffer_755 = _RAND_755[15:0];
  _RAND_756 = {1{`RANDOM}};
  buffer_756 = _RAND_756[15:0];
  _RAND_757 = {1{`RANDOM}};
  buffer_757 = _RAND_757[15:0];
  _RAND_758 = {1{`RANDOM}};
  buffer_758 = _RAND_758[15:0];
  _RAND_759 = {1{`RANDOM}};
  buffer_759 = _RAND_759[15:0];
  _RAND_760 = {1{`RANDOM}};
  buffer_760 = _RAND_760[15:0];
  _RAND_761 = {1{`RANDOM}};
  buffer_761 = _RAND_761[15:0];
  _RAND_762 = {1{`RANDOM}};
  buffer_762 = _RAND_762[15:0];
  _RAND_763 = {1{`RANDOM}};
  buffer_763 = _RAND_763[15:0];
  _RAND_764 = {1{`RANDOM}};
  buffer_764 = _RAND_764[15:0];
  _RAND_765 = {1{`RANDOM}};
  buffer_765 = _RAND_765[15:0];
  _RAND_766 = {1{`RANDOM}};
  buffer_766 = _RAND_766[15:0];
  _RAND_767 = {1{`RANDOM}};
  buffer_767 = _RAND_767[15:0];
  _RAND_768 = {1{`RANDOM}};
  buffer_768 = _RAND_768[15:0];
  _RAND_769 = {1{`RANDOM}};
  buffer_769 = _RAND_769[15:0];
  _RAND_770 = {1{`RANDOM}};
  buffer_770 = _RAND_770[15:0];
  _RAND_771 = {1{`RANDOM}};
  buffer_771 = _RAND_771[15:0];
  _RAND_772 = {1{`RANDOM}};
  buffer_772 = _RAND_772[15:0];
  _RAND_773 = {1{`RANDOM}};
  buffer_773 = _RAND_773[15:0];
  _RAND_774 = {1{`RANDOM}};
  buffer_774 = _RAND_774[15:0];
  _RAND_775 = {1{`RANDOM}};
  buffer_775 = _RAND_775[15:0];
  _RAND_776 = {1{`RANDOM}};
  buffer_776 = _RAND_776[15:0];
  _RAND_777 = {1{`RANDOM}};
  buffer_777 = _RAND_777[15:0];
  _RAND_778 = {1{`RANDOM}};
  buffer_778 = _RAND_778[15:0];
  _RAND_779 = {1{`RANDOM}};
  buffer_779 = _RAND_779[15:0];
  _RAND_780 = {1{`RANDOM}};
  buffer_780 = _RAND_780[15:0];
  _RAND_781 = {1{`RANDOM}};
  buffer_781 = _RAND_781[15:0];
  _RAND_782 = {1{`RANDOM}};
  buffer_782 = _RAND_782[15:0];
  _RAND_783 = {1{`RANDOM}};
  buffer_783 = _RAND_783[15:0];
  _RAND_784 = {1{`RANDOM}};
  buffer_784 = _RAND_784[15:0];
  _RAND_785 = {1{`RANDOM}};
  buffer_785 = _RAND_785[15:0];
  _RAND_786 = {1{`RANDOM}};
  buffer_786 = _RAND_786[15:0];
  _RAND_787 = {1{`RANDOM}};
  buffer_787 = _RAND_787[15:0];
  _RAND_788 = {1{`RANDOM}};
  buffer_788 = _RAND_788[15:0];
  _RAND_789 = {1{`RANDOM}};
  buffer_789 = _RAND_789[15:0];
  _RAND_790 = {1{`RANDOM}};
  buffer_790 = _RAND_790[15:0];
  _RAND_791 = {1{`RANDOM}};
  buffer_791 = _RAND_791[15:0];
  _RAND_792 = {1{`RANDOM}};
  buffer_792 = _RAND_792[15:0];
  _RAND_793 = {1{`RANDOM}};
  buffer_793 = _RAND_793[15:0];
  _RAND_794 = {1{`RANDOM}};
  buffer_794 = _RAND_794[15:0];
  _RAND_795 = {1{`RANDOM}};
  buffer_795 = _RAND_795[15:0];
  _RAND_796 = {1{`RANDOM}};
  buffer_796 = _RAND_796[15:0];
  _RAND_797 = {1{`RANDOM}};
  buffer_797 = _RAND_797[15:0];
  _RAND_798 = {1{`RANDOM}};
  buffer_798 = _RAND_798[15:0];
  _RAND_799 = {1{`RANDOM}};
  buffer_799 = _RAND_799[15:0];
  _RAND_800 = {1{`RANDOM}};
  buffer_800 = _RAND_800[15:0];
  _RAND_801 = {1{`RANDOM}};
  buffer_801 = _RAND_801[15:0];
  _RAND_802 = {1{`RANDOM}};
  buffer_802 = _RAND_802[15:0];
  _RAND_803 = {1{`RANDOM}};
  buffer_803 = _RAND_803[15:0];
  _RAND_804 = {1{`RANDOM}};
  buffer_804 = _RAND_804[15:0];
  _RAND_805 = {1{`RANDOM}};
  buffer_805 = _RAND_805[15:0];
  _RAND_806 = {1{`RANDOM}};
  buffer_806 = _RAND_806[15:0];
  _RAND_807 = {1{`RANDOM}};
  buffer_807 = _RAND_807[15:0];
  _RAND_808 = {1{`RANDOM}};
  buffer_808 = _RAND_808[15:0];
  _RAND_809 = {1{`RANDOM}};
  buffer_809 = _RAND_809[15:0];
  _RAND_810 = {1{`RANDOM}};
  buffer_810 = _RAND_810[15:0];
  _RAND_811 = {1{`RANDOM}};
  buffer_811 = _RAND_811[15:0];
  _RAND_812 = {1{`RANDOM}};
  buffer_812 = _RAND_812[15:0];
  _RAND_813 = {1{`RANDOM}};
  buffer_813 = _RAND_813[15:0];
  _RAND_814 = {1{`RANDOM}};
  buffer_814 = _RAND_814[15:0];
  _RAND_815 = {1{`RANDOM}};
  buffer_815 = _RAND_815[15:0];
  _RAND_816 = {1{`RANDOM}};
  buffer_816 = _RAND_816[15:0];
  _RAND_817 = {1{`RANDOM}};
  buffer_817 = _RAND_817[15:0];
  _RAND_818 = {1{`RANDOM}};
  buffer_818 = _RAND_818[15:0];
  _RAND_819 = {1{`RANDOM}};
  buffer_819 = _RAND_819[15:0];
  _RAND_820 = {1{`RANDOM}};
  buffer_820 = _RAND_820[15:0];
  _RAND_821 = {1{`RANDOM}};
  buffer_821 = _RAND_821[15:0];
  _RAND_822 = {1{`RANDOM}};
  buffer_822 = _RAND_822[15:0];
  _RAND_823 = {1{`RANDOM}};
  buffer_823 = _RAND_823[15:0];
  _RAND_824 = {1{`RANDOM}};
  buffer_824 = _RAND_824[15:0];
  _RAND_825 = {1{`RANDOM}};
  buffer_825 = _RAND_825[15:0];
  _RAND_826 = {1{`RANDOM}};
  buffer_826 = _RAND_826[15:0];
  _RAND_827 = {1{`RANDOM}};
  buffer_827 = _RAND_827[15:0];
  _RAND_828 = {1{`RANDOM}};
  buffer_828 = _RAND_828[15:0];
  _RAND_829 = {1{`RANDOM}};
  buffer_829 = _RAND_829[15:0];
  _RAND_830 = {1{`RANDOM}};
  buffer_830 = _RAND_830[15:0];
  _RAND_831 = {1{`RANDOM}};
  buffer_831 = _RAND_831[15:0];
  _RAND_832 = {1{`RANDOM}};
  buffer_832 = _RAND_832[15:0];
  _RAND_833 = {1{`RANDOM}};
  buffer_833 = _RAND_833[15:0];
  _RAND_834 = {1{`RANDOM}};
  buffer_834 = _RAND_834[15:0];
  _RAND_835 = {1{`RANDOM}};
  buffer_835 = _RAND_835[15:0];
  _RAND_836 = {1{`RANDOM}};
  buffer_836 = _RAND_836[15:0];
  _RAND_837 = {1{`RANDOM}};
  buffer_837 = _RAND_837[15:0];
  _RAND_838 = {1{`RANDOM}};
  buffer_838 = _RAND_838[15:0];
  _RAND_839 = {1{`RANDOM}};
  buffer_839 = _RAND_839[15:0];
  _RAND_840 = {1{`RANDOM}};
  buffer_840 = _RAND_840[15:0];
  _RAND_841 = {1{`RANDOM}};
  buffer_841 = _RAND_841[15:0];
  _RAND_842 = {1{`RANDOM}};
  buffer_842 = _RAND_842[15:0];
  _RAND_843 = {1{`RANDOM}};
  buffer_843 = _RAND_843[15:0];
  _RAND_844 = {1{`RANDOM}};
  buffer_844 = _RAND_844[15:0];
  _RAND_845 = {1{`RANDOM}};
  buffer_845 = _RAND_845[15:0];
  _RAND_846 = {1{`RANDOM}};
  buffer_846 = _RAND_846[15:0];
  _RAND_847 = {1{`RANDOM}};
  buffer_847 = _RAND_847[15:0];
  _RAND_848 = {1{`RANDOM}};
  buffer_848 = _RAND_848[15:0];
  _RAND_849 = {1{`RANDOM}};
  buffer_849 = _RAND_849[15:0];
  _RAND_850 = {1{`RANDOM}};
  buffer_850 = _RAND_850[15:0];
  _RAND_851 = {1{`RANDOM}};
  buffer_851 = _RAND_851[15:0];
  _RAND_852 = {1{`RANDOM}};
  buffer_852 = _RAND_852[15:0];
  _RAND_853 = {1{`RANDOM}};
  buffer_853 = _RAND_853[15:0];
  _RAND_854 = {1{`RANDOM}};
  buffer_854 = _RAND_854[15:0];
  _RAND_855 = {1{`RANDOM}};
  buffer_855 = _RAND_855[15:0];
  _RAND_856 = {1{`RANDOM}};
  buffer_856 = _RAND_856[15:0];
  _RAND_857 = {1{`RANDOM}};
  buffer_857 = _RAND_857[15:0];
  _RAND_858 = {1{`RANDOM}};
  buffer_858 = _RAND_858[15:0];
  _RAND_859 = {1{`RANDOM}};
  buffer_859 = _RAND_859[15:0];
  _RAND_860 = {1{`RANDOM}};
  buffer_860 = _RAND_860[15:0];
  _RAND_861 = {1{`RANDOM}};
  buffer_861 = _RAND_861[15:0];
  _RAND_862 = {1{`RANDOM}};
  buffer_862 = _RAND_862[15:0];
  _RAND_863 = {1{`RANDOM}};
  buffer_863 = _RAND_863[15:0];
  _RAND_864 = {1{`RANDOM}};
  buffer_864 = _RAND_864[15:0];
  _RAND_865 = {1{`RANDOM}};
  buffer_865 = _RAND_865[15:0];
  _RAND_866 = {1{`RANDOM}};
  buffer_866 = _RAND_866[15:0];
  _RAND_867 = {1{`RANDOM}};
  buffer_867 = _RAND_867[15:0];
  _RAND_868 = {1{`RANDOM}};
  buffer_868 = _RAND_868[15:0];
  _RAND_869 = {1{`RANDOM}};
  buffer_869 = _RAND_869[15:0];
  _RAND_870 = {1{`RANDOM}};
  buffer_870 = _RAND_870[15:0];
  _RAND_871 = {1{`RANDOM}};
  buffer_871 = _RAND_871[15:0];
  _RAND_872 = {1{`RANDOM}};
  buffer_872 = _RAND_872[15:0];
  _RAND_873 = {1{`RANDOM}};
  buffer_873 = _RAND_873[15:0];
  _RAND_874 = {1{`RANDOM}};
  buffer_874 = _RAND_874[15:0];
  _RAND_875 = {1{`RANDOM}};
  buffer_875 = _RAND_875[15:0];
  _RAND_876 = {1{`RANDOM}};
  buffer_876 = _RAND_876[15:0];
  _RAND_877 = {1{`RANDOM}};
  buffer_877 = _RAND_877[15:0];
  _RAND_878 = {1{`RANDOM}};
  buffer_878 = _RAND_878[15:0];
  _RAND_879 = {1{`RANDOM}};
  buffer_879 = _RAND_879[15:0];
  _RAND_880 = {1{`RANDOM}};
  buffer_880 = _RAND_880[15:0];
  _RAND_881 = {1{`RANDOM}};
  buffer_881 = _RAND_881[15:0];
  _RAND_882 = {1{`RANDOM}};
  buffer_882 = _RAND_882[15:0];
  _RAND_883 = {1{`RANDOM}};
  buffer_883 = _RAND_883[15:0];
  _RAND_884 = {1{`RANDOM}};
  buffer_884 = _RAND_884[15:0];
  _RAND_885 = {1{`RANDOM}};
  buffer_885 = _RAND_885[15:0];
  _RAND_886 = {1{`RANDOM}};
  buffer_886 = _RAND_886[15:0];
  _RAND_887 = {1{`RANDOM}};
  buffer_887 = _RAND_887[15:0];
  _RAND_888 = {1{`RANDOM}};
  buffer_888 = _RAND_888[15:0];
  _RAND_889 = {1{`RANDOM}};
  buffer_889 = _RAND_889[15:0];
  _RAND_890 = {1{`RANDOM}};
  buffer_890 = _RAND_890[15:0];
  _RAND_891 = {1{`RANDOM}};
  buffer_891 = _RAND_891[15:0];
  _RAND_892 = {1{`RANDOM}};
  buffer_892 = _RAND_892[15:0];
  _RAND_893 = {1{`RANDOM}};
  buffer_893 = _RAND_893[15:0];
  _RAND_894 = {1{`RANDOM}};
  buffer_894 = _RAND_894[15:0];
  _RAND_895 = {1{`RANDOM}};
  buffer_895 = _RAND_895[15:0];
  _RAND_896 = {1{`RANDOM}};
  buffer_896 = _RAND_896[15:0];
  _RAND_897 = {1{`RANDOM}};
  buffer_897 = _RAND_897[15:0];
  _RAND_898 = {1{`RANDOM}};
  buffer_898 = _RAND_898[15:0];
  _RAND_899 = {1{`RANDOM}};
  buffer_899 = _RAND_899[15:0];
  _RAND_900 = {1{`RANDOM}};
  buffer_900 = _RAND_900[15:0];
  _RAND_901 = {1{`RANDOM}};
  buffer_901 = _RAND_901[15:0];
  _RAND_902 = {1{`RANDOM}};
  buffer_902 = _RAND_902[15:0];
  _RAND_903 = {1{`RANDOM}};
  buffer_903 = _RAND_903[15:0];
  _RAND_904 = {1{`RANDOM}};
  buffer_904 = _RAND_904[15:0];
  _RAND_905 = {1{`RANDOM}};
  buffer_905 = _RAND_905[15:0];
  _RAND_906 = {1{`RANDOM}};
  buffer_906 = _RAND_906[15:0];
  _RAND_907 = {1{`RANDOM}};
  buffer_907 = _RAND_907[15:0];
  _RAND_908 = {1{`RANDOM}};
  buffer_908 = _RAND_908[15:0];
  _RAND_909 = {1{`RANDOM}};
  buffer_909 = _RAND_909[15:0];
  _RAND_910 = {1{`RANDOM}};
  buffer_910 = _RAND_910[15:0];
  _RAND_911 = {1{`RANDOM}};
  buffer_911 = _RAND_911[15:0];
  _RAND_912 = {1{`RANDOM}};
  buffer_912 = _RAND_912[15:0];
  _RAND_913 = {1{`RANDOM}};
  buffer_913 = _RAND_913[15:0];
  _RAND_914 = {1{`RANDOM}};
  buffer_914 = _RAND_914[15:0];
  _RAND_915 = {1{`RANDOM}};
  buffer_915 = _RAND_915[15:0];
  _RAND_916 = {1{`RANDOM}};
  buffer_916 = _RAND_916[15:0];
  _RAND_917 = {1{`RANDOM}};
  buffer_917 = _RAND_917[15:0];
  _RAND_918 = {1{`RANDOM}};
  buffer_918 = _RAND_918[15:0];
  _RAND_919 = {1{`RANDOM}};
  buffer_919 = _RAND_919[15:0];
  _RAND_920 = {1{`RANDOM}};
  buffer_920 = _RAND_920[15:0];
  _RAND_921 = {1{`RANDOM}};
  buffer_921 = _RAND_921[15:0];
  _RAND_922 = {1{`RANDOM}};
  buffer_922 = _RAND_922[15:0];
  _RAND_923 = {1{`RANDOM}};
  buffer_923 = _RAND_923[15:0];
  _RAND_924 = {1{`RANDOM}};
  buffer_924 = _RAND_924[15:0];
  _RAND_925 = {1{`RANDOM}};
  buffer_925 = _RAND_925[15:0];
  _RAND_926 = {1{`RANDOM}};
  buffer_926 = _RAND_926[15:0];
  _RAND_927 = {1{`RANDOM}};
  buffer_927 = _RAND_927[15:0];
  _RAND_928 = {1{`RANDOM}};
  buffer_928 = _RAND_928[15:0];
  _RAND_929 = {1{`RANDOM}};
  buffer_929 = _RAND_929[15:0];
  _RAND_930 = {1{`RANDOM}};
  buffer_930 = _RAND_930[15:0];
  _RAND_931 = {1{`RANDOM}};
  buffer_931 = _RAND_931[15:0];
  _RAND_932 = {1{`RANDOM}};
  buffer_932 = _RAND_932[15:0];
  _RAND_933 = {1{`RANDOM}};
  buffer_933 = _RAND_933[15:0];
  _RAND_934 = {1{`RANDOM}};
  buffer_934 = _RAND_934[15:0];
  _RAND_935 = {1{`RANDOM}};
  buffer_935 = _RAND_935[15:0];
  _RAND_936 = {1{`RANDOM}};
  buffer_936 = _RAND_936[15:0];
  _RAND_937 = {1{`RANDOM}};
  buffer_937 = _RAND_937[15:0];
  _RAND_938 = {1{`RANDOM}};
  buffer_938 = _RAND_938[15:0];
  _RAND_939 = {1{`RANDOM}};
  buffer_939 = _RAND_939[15:0];
  _RAND_940 = {1{`RANDOM}};
  buffer_940 = _RAND_940[15:0];
  _RAND_941 = {1{`RANDOM}};
  buffer_941 = _RAND_941[15:0];
  _RAND_942 = {1{`RANDOM}};
  buffer_942 = _RAND_942[15:0];
  _RAND_943 = {1{`RANDOM}};
  buffer_943 = _RAND_943[15:0];
  _RAND_944 = {1{`RANDOM}};
  buffer_944 = _RAND_944[15:0];
  _RAND_945 = {1{`RANDOM}};
  buffer_945 = _RAND_945[15:0];
  _RAND_946 = {1{`RANDOM}};
  buffer_946 = _RAND_946[15:0];
  _RAND_947 = {1{`RANDOM}};
  buffer_947 = _RAND_947[15:0];
  _RAND_948 = {1{`RANDOM}};
  buffer_948 = _RAND_948[15:0];
  _RAND_949 = {1{`RANDOM}};
  buffer_949 = _RAND_949[15:0];
  _RAND_950 = {1{`RANDOM}};
  buffer_950 = _RAND_950[15:0];
  _RAND_951 = {1{`RANDOM}};
  buffer_951 = _RAND_951[15:0];
  _RAND_952 = {1{`RANDOM}};
  buffer_952 = _RAND_952[15:0];
  _RAND_953 = {1{`RANDOM}};
  buffer_953 = _RAND_953[15:0];
  _RAND_954 = {1{`RANDOM}};
  buffer_954 = _RAND_954[15:0];
  _RAND_955 = {1{`RANDOM}};
  buffer_955 = _RAND_955[15:0];
  _RAND_956 = {1{`RANDOM}};
  buffer_956 = _RAND_956[15:0];
  _RAND_957 = {1{`RANDOM}};
  buffer_957 = _RAND_957[15:0];
  _RAND_958 = {1{`RANDOM}};
  buffer_958 = _RAND_958[15:0];
  _RAND_959 = {1{`RANDOM}};
  buffer_959 = _RAND_959[15:0];
  _RAND_960 = {1{`RANDOM}};
  buffer_960 = _RAND_960[15:0];
  _RAND_961 = {1{`RANDOM}};
  buffer_961 = _RAND_961[15:0];
  _RAND_962 = {1{`RANDOM}};
  buffer_962 = _RAND_962[15:0];
  _RAND_963 = {1{`RANDOM}};
  buffer_963 = _RAND_963[15:0];
  _RAND_964 = {1{`RANDOM}};
  buffer_964 = _RAND_964[15:0];
  _RAND_965 = {1{`RANDOM}};
  buffer_965 = _RAND_965[15:0];
  _RAND_966 = {1{`RANDOM}};
  buffer_966 = _RAND_966[15:0];
  _RAND_967 = {1{`RANDOM}};
  buffer_967 = _RAND_967[15:0];
  _RAND_968 = {1{`RANDOM}};
  buffer_968 = _RAND_968[15:0];
  _RAND_969 = {1{`RANDOM}};
  buffer_969 = _RAND_969[15:0];
  _RAND_970 = {1{`RANDOM}};
  buffer_970 = _RAND_970[15:0];
  _RAND_971 = {1{`RANDOM}};
  buffer_971 = _RAND_971[15:0];
  _RAND_972 = {1{`RANDOM}};
  buffer_972 = _RAND_972[15:0];
  _RAND_973 = {1{`RANDOM}};
  buffer_973 = _RAND_973[15:0];
  _RAND_974 = {1{`RANDOM}};
  buffer_974 = _RAND_974[15:0];
  _RAND_975 = {1{`RANDOM}};
  buffer_975 = _RAND_975[15:0];
  _RAND_976 = {1{`RANDOM}};
  buffer_976 = _RAND_976[15:0];
  _RAND_977 = {1{`RANDOM}};
  buffer_977 = _RAND_977[15:0];
  _RAND_978 = {1{`RANDOM}};
  buffer_978 = _RAND_978[15:0];
  _RAND_979 = {1{`RANDOM}};
  buffer_979 = _RAND_979[15:0];
  _RAND_980 = {1{`RANDOM}};
  buffer_980 = _RAND_980[15:0];
  _RAND_981 = {1{`RANDOM}};
  buffer_981 = _RAND_981[15:0];
  _RAND_982 = {1{`RANDOM}};
  buffer_982 = _RAND_982[15:0];
  _RAND_983 = {1{`RANDOM}};
  buffer_983 = _RAND_983[15:0];
  _RAND_984 = {1{`RANDOM}};
  buffer_984 = _RAND_984[15:0];
  _RAND_985 = {1{`RANDOM}};
  buffer_985 = _RAND_985[15:0];
  _RAND_986 = {1{`RANDOM}};
  buffer_986 = _RAND_986[15:0];
  _RAND_987 = {1{`RANDOM}};
  buffer_987 = _RAND_987[15:0];
  _RAND_988 = {1{`RANDOM}};
  buffer_988 = _RAND_988[15:0];
  _RAND_989 = {1{`RANDOM}};
  buffer_989 = _RAND_989[15:0];
  _RAND_990 = {1{`RANDOM}};
  buffer_990 = _RAND_990[15:0];
  _RAND_991 = {1{`RANDOM}};
  buffer_991 = _RAND_991[15:0];
  _RAND_992 = {1{`RANDOM}};
  buffer_992 = _RAND_992[15:0];
  _RAND_993 = {1{`RANDOM}};
  buffer_993 = _RAND_993[15:0];
  _RAND_994 = {1{`RANDOM}};
  buffer_994 = _RAND_994[15:0];
  _RAND_995 = {1{`RANDOM}};
  buffer_995 = _RAND_995[15:0];
  _RAND_996 = {1{`RANDOM}};
  buffer_996 = _RAND_996[15:0];
  _RAND_997 = {1{`RANDOM}};
  buffer_997 = _RAND_997[15:0];
  _RAND_998 = {1{`RANDOM}};
  buffer_998 = _RAND_998[15:0];
  _RAND_999 = {1{`RANDOM}};
  buffer_999 = _RAND_999[15:0];
  _RAND_1000 = {1{`RANDOM}};
  buffer_1000 = _RAND_1000[15:0];
  _RAND_1001 = {1{`RANDOM}};
  buffer_1001 = _RAND_1001[15:0];
  _RAND_1002 = {1{`RANDOM}};
  buffer_1002 = _RAND_1002[15:0];
  _RAND_1003 = {1{`RANDOM}};
  buffer_1003 = _RAND_1003[15:0];
  _RAND_1004 = {1{`RANDOM}};
  buffer_1004 = _RAND_1004[15:0];
  _RAND_1005 = {1{`RANDOM}};
  buffer_1005 = _RAND_1005[15:0];
  _RAND_1006 = {1{`RANDOM}};
  buffer_1006 = _RAND_1006[15:0];
  _RAND_1007 = {1{`RANDOM}};
  buffer_1007 = _RAND_1007[15:0];
  _RAND_1008 = {1{`RANDOM}};
  buffer_1008 = _RAND_1008[15:0];
  _RAND_1009 = {1{`RANDOM}};
  buffer_1009 = _RAND_1009[15:0];
  _RAND_1010 = {1{`RANDOM}};
  buffer_1010 = _RAND_1010[15:0];
  _RAND_1011 = {1{`RANDOM}};
  buffer_1011 = _RAND_1011[15:0];
  _RAND_1012 = {1{`RANDOM}};
  buffer_1012 = _RAND_1012[15:0];
  _RAND_1013 = {1{`RANDOM}};
  buffer_1013 = _RAND_1013[15:0];
  _RAND_1014 = {1{`RANDOM}};
  buffer_1014 = _RAND_1014[15:0];
  _RAND_1015 = {1{`RANDOM}};
  buffer_1015 = _RAND_1015[15:0];
  _RAND_1016 = {1{`RANDOM}};
  buffer_1016 = _RAND_1016[15:0];
  _RAND_1017 = {1{`RANDOM}};
  buffer_1017 = _RAND_1017[15:0];
  _RAND_1018 = {1{`RANDOM}};
  buffer_1018 = _RAND_1018[15:0];
  _RAND_1019 = {1{`RANDOM}};
  buffer_1019 = _RAND_1019[15:0];
  _RAND_1020 = {1{`RANDOM}};
  buffer_1020 = _RAND_1020[15:0];
  _RAND_1021 = {1{`RANDOM}};
  buffer_1021 = _RAND_1021[15:0];
  _RAND_1022 = {1{`RANDOM}};
  buffer_1022 = _RAND_1022[15:0];
  _RAND_1023 = {1{`RANDOM}};
  buffer_1023 = _RAND_1023[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module OuterBuffer(
  input         clock,
  input         reset,
  input  [15:0] io_BufferIO_DataIn,
  input  [9:0]  io_BufferIO_DataAddr,
  input         io_BufferIO_ReadWrite,
  input         io_BufferIO_Enable,
  output [15:0] io_BufferIO_DataOut,
  input  [3:0]  io_BankIndex
);
  wire  bank0_clock; // @[OuterBuffer.scala 41:23]
  wire  bank0_reset; // @[OuterBuffer.scala 41:23]
  wire [15:0] bank0_io_BankIO_DataIn; // @[OuterBuffer.scala 41:23]
  wire [9:0] bank0_io_BankIO_DataAddr; // @[OuterBuffer.scala 41:23]
  wire  bank0_io_BankIO_ReadWrite; // @[OuterBuffer.scala 41:23]
  wire  bank0_io_BankIO_Enable; // @[OuterBuffer.scala 41:23]
  wire [15:0] bank0_io_BankIO_DataOut; // @[OuterBuffer.scala 41:23]
  wire  bank1_clock; // @[OuterBuffer.scala 42:23]
  wire  bank1_reset; // @[OuterBuffer.scala 42:23]
  wire [15:0] bank1_io_BankIO_DataIn; // @[OuterBuffer.scala 42:23]
  wire [9:0] bank1_io_BankIO_DataAddr; // @[OuterBuffer.scala 42:23]
  wire  bank1_io_BankIO_ReadWrite; // @[OuterBuffer.scala 42:23]
  wire  bank1_io_BankIO_Enable; // @[OuterBuffer.scala 42:23]
  wire [15:0] bank1_io_BankIO_DataOut; // @[OuterBuffer.scala 42:23]
  wire  bank2_clock; // @[OuterBuffer.scala 43:23]
  wire  bank2_reset; // @[OuterBuffer.scala 43:23]
  wire [15:0] bank2_io_BankIO_DataIn; // @[OuterBuffer.scala 43:23]
  wire [9:0] bank2_io_BankIO_DataAddr; // @[OuterBuffer.scala 43:23]
  wire  bank2_io_BankIO_ReadWrite; // @[OuterBuffer.scala 43:23]
  wire  bank2_io_BankIO_Enable; // @[OuterBuffer.scala 43:23]
  wire [15:0] bank2_io_BankIO_DataOut; // @[OuterBuffer.scala 43:23]
  wire  bank3_clock; // @[OuterBuffer.scala 44:23]
  wire  bank3_reset; // @[OuterBuffer.scala 44:23]
  wire [15:0] bank3_io_BankIO_DataIn; // @[OuterBuffer.scala 44:23]
  wire [9:0] bank3_io_BankIO_DataAddr; // @[OuterBuffer.scala 44:23]
  wire  bank3_io_BankIO_ReadWrite; // @[OuterBuffer.scala 44:23]
  wire  bank3_io_BankIO_Enable; // @[OuterBuffer.scala 44:23]
  wire [15:0] bank3_io_BankIO_DataOut; // @[OuterBuffer.scala 44:23]
  wire  bank4_clock; // @[OuterBuffer.scala 45:23]
  wire  bank4_reset; // @[OuterBuffer.scala 45:23]
  wire [15:0] bank4_io_BankIO_DataIn; // @[OuterBuffer.scala 45:23]
  wire [9:0] bank4_io_BankIO_DataAddr; // @[OuterBuffer.scala 45:23]
  wire  bank4_io_BankIO_ReadWrite; // @[OuterBuffer.scala 45:23]
  wire  bank4_io_BankIO_Enable; // @[OuterBuffer.scala 45:23]
  wire [15:0] bank4_io_BankIO_DataOut; // @[OuterBuffer.scala 45:23]
  wire  bank5_clock; // @[OuterBuffer.scala 46:23]
  wire  bank5_reset; // @[OuterBuffer.scala 46:23]
  wire [15:0] bank5_io_BankIO_DataIn; // @[OuterBuffer.scala 46:23]
  wire [9:0] bank5_io_BankIO_DataAddr; // @[OuterBuffer.scala 46:23]
  wire  bank5_io_BankIO_ReadWrite; // @[OuterBuffer.scala 46:23]
  wire  bank5_io_BankIO_Enable; // @[OuterBuffer.scala 46:23]
  wire [15:0] bank5_io_BankIO_DataOut; // @[OuterBuffer.scala 46:23]
  wire  bank6_clock; // @[OuterBuffer.scala 47:23]
  wire  bank6_reset; // @[OuterBuffer.scala 47:23]
  wire [15:0] bank6_io_BankIO_DataIn; // @[OuterBuffer.scala 47:23]
  wire [9:0] bank6_io_BankIO_DataAddr; // @[OuterBuffer.scala 47:23]
  wire  bank6_io_BankIO_ReadWrite; // @[OuterBuffer.scala 47:23]
  wire  bank6_io_BankIO_Enable; // @[OuterBuffer.scala 47:23]
  wire [15:0] bank6_io_BankIO_DataOut; // @[OuterBuffer.scala 47:23]
  wire  bank7_clock; // @[OuterBuffer.scala 48:23]
  wire  bank7_reset; // @[OuterBuffer.scala 48:23]
  wire [15:0] bank7_io_BankIO_DataIn; // @[OuterBuffer.scala 48:23]
  wire [9:0] bank7_io_BankIO_DataAddr; // @[OuterBuffer.scala 48:23]
  wire  bank7_io_BankIO_ReadWrite; // @[OuterBuffer.scala 48:23]
  wire  bank7_io_BankIO_Enable; // @[OuterBuffer.scala 48:23]
  wire [15:0] bank7_io_BankIO_DataOut; // @[OuterBuffer.scala 48:23]
  wire  bank8_clock; // @[OuterBuffer.scala 49:23]
  wire  bank8_reset; // @[OuterBuffer.scala 49:23]
  wire [15:0] bank8_io_BankIO_DataIn; // @[OuterBuffer.scala 49:23]
  wire [9:0] bank8_io_BankIO_DataAddr; // @[OuterBuffer.scala 49:23]
  wire  bank8_io_BankIO_ReadWrite; // @[OuterBuffer.scala 49:23]
  wire  bank8_io_BankIO_Enable; // @[OuterBuffer.scala 49:23]
  wire [15:0] bank8_io_BankIO_DataOut; // @[OuterBuffer.scala 49:23]
  wire  bank9_clock; // @[OuterBuffer.scala 50:23]
  wire  bank9_reset; // @[OuterBuffer.scala 50:23]
  wire [15:0] bank9_io_BankIO_DataIn; // @[OuterBuffer.scala 50:23]
  wire [9:0] bank9_io_BankIO_DataAddr; // @[OuterBuffer.scala 50:23]
  wire  bank9_io_BankIO_ReadWrite; // @[OuterBuffer.scala 50:23]
  wire  bank9_io_BankIO_Enable; // @[OuterBuffer.scala 50:23]
  wire [15:0] bank9_io_BankIO_DataOut; // @[OuterBuffer.scala 50:23]
  wire  bank10_clock; // @[OuterBuffer.scala 51:23]
  wire  bank10_reset; // @[OuterBuffer.scala 51:23]
  wire [15:0] bank10_io_BankIO_DataIn; // @[OuterBuffer.scala 51:23]
  wire [9:0] bank10_io_BankIO_DataAddr; // @[OuterBuffer.scala 51:23]
  wire  bank10_io_BankIO_ReadWrite; // @[OuterBuffer.scala 51:23]
  wire  bank10_io_BankIO_Enable; // @[OuterBuffer.scala 51:23]
  wire [15:0] bank10_io_BankIO_DataOut; // @[OuterBuffer.scala 51:23]
  wire  bank11_clock; // @[OuterBuffer.scala 52:23]
  wire  bank11_reset; // @[OuterBuffer.scala 52:23]
  wire [15:0] bank11_io_BankIO_DataIn; // @[OuterBuffer.scala 52:23]
  wire [9:0] bank11_io_BankIO_DataAddr; // @[OuterBuffer.scala 52:23]
  wire  bank11_io_BankIO_ReadWrite; // @[OuterBuffer.scala 52:23]
  wire  bank11_io_BankIO_Enable; // @[OuterBuffer.scala 52:23]
  wire [15:0] bank11_io_BankIO_DataOut; // @[OuterBuffer.scala 52:23]
  wire  bank12_clock; // @[OuterBuffer.scala 53:23]
  wire  bank12_reset; // @[OuterBuffer.scala 53:23]
  wire [15:0] bank12_io_BankIO_DataIn; // @[OuterBuffer.scala 53:23]
  wire [9:0] bank12_io_BankIO_DataAddr; // @[OuterBuffer.scala 53:23]
  wire  bank12_io_BankIO_ReadWrite; // @[OuterBuffer.scala 53:23]
  wire  bank12_io_BankIO_Enable; // @[OuterBuffer.scala 53:23]
  wire [15:0] bank12_io_BankIO_DataOut; // @[OuterBuffer.scala 53:23]
  wire  bank13_clock; // @[OuterBuffer.scala 54:23]
  wire  bank13_reset; // @[OuterBuffer.scala 54:23]
  wire [15:0] bank13_io_BankIO_DataIn; // @[OuterBuffer.scala 54:23]
  wire [9:0] bank13_io_BankIO_DataAddr; // @[OuterBuffer.scala 54:23]
  wire  bank13_io_BankIO_ReadWrite; // @[OuterBuffer.scala 54:23]
  wire  bank13_io_BankIO_Enable; // @[OuterBuffer.scala 54:23]
  wire [15:0] bank13_io_BankIO_DataOut; // @[OuterBuffer.scala 54:23]
  wire  bank14_clock; // @[OuterBuffer.scala 55:23]
  wire  bank14_reset; // @[OuterBuffer.scala 55:23]
  wire [15:0] bank14_io_BankIO_DataIn; // @[OuterBuffer.scala 55:23]
  wire [9:0] bank14_io_BankIO_DataAddr; // @[OuterBuffer.scala 55:23]
  wire  bank14_io_BankIO_ReadWrite; // @[OuterBuffer.scala 55:23]
  wire  bank14_io_BankIO_Enable; // @[OuterBuffer.scala 55:23]
  wire [15:0] bank14_io_BankIO_DataOut; // @[OuterBuffer.scala 55:23]
  wire  bank15_clock; // @[OuterBuffer.scala 56:23]
  wire  bank15_reset; // @[OuterBuffer.scala 56:23]
  wire [15:0] bank15_io_BankIO_DataIn; // @[OuterBuffer.scala 56:23]
  wire [9:0] bank15_io_BankIO_DataAddr; // @[OuterBuffer.scala 56:23]
  wire  bank15_io_BankIO_ReadWrite; // @[OuterBuffer.scala 56:23]
  wire  bank15_io_BankIO_Enable; // @[OuterBuffer.scala 56:23]
  wire [15:0] bank15_io_BankIO_DataOut; // @[OuterBuffer.scala 56:23]
  wire  _T = 4'h0 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_1 = 4'h1 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_2 = 4'h2 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_3 = 4'h3 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_4 = 4'h4 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_5 = 4'h5 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_6 = 4'h6 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_7 = 4'h7 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_8 = 4'h8 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_9 = 4'h9 == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_10 = 4'ha == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_11 = 4'hb == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_12 = 4'hc == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_13 = 4'hd == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_14 = 4'he == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _T_15 = 4'hf == io_BankIndex; // @[OuterBuffer.scala 95:24]
  wire  _GEN_0 = 4'hf == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 111:40 91:27]
  wire  _GEN_1 = 4'he == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 110:40 90:27]
  wire  _GEN_2 = 4'he == io_BankIndex ? 1'h0 : _GEN_0; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_3 = 4'hd == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 109:40 89:27]
  wire  _GEN_4 = 4'hd == io_BankIndex ? 1'h0 : _GEN_1; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_5 = 4'hd == io_BankIndex ? 1'h0 : _GEN_2; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_6 = 4'hc == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 108:40 88:27]
  wire  _GEN_7 = 4'hc == io_BankIndex ? 1'h0 : _GEN_3; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_8 = 4'hc == io_BankIndex ? 1'h0 : _GEN_4; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_9 = 4'hc == io_BankIndex ? 1'h0 : _GEN_5; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_10 = 4'hb == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 107:40 87:27]
  wire  _GEN_11 = 4'hb == io_BankIndex ? 1'h0 : _GEN_6; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_12 = 4'hb == io_BankIndex ? 1'h0 : _GEN_7; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_13 = 4'hb == io_BankIndex ? 1'h0 : _GEN_8; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_14 = 4'hb == io_BankIndex ? 1'h0 : _GEN_9; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_15 = 4'ha == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 106:40 86:27]
  wire  _GEN_16 = 4'ha == io_BankIndex ? 1'h0 : _GEN_10; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_17 = 4'ha == io_BankIndex ? 1'h0 : _GEN_11; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_18 = 4'ha == io_BankIndex ? 1'h0 : _GEN_12; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_19 = 4'ha == io_BankIndex ? 1'h0 : _GEN_13; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_20 = 4'ha == io_BankIndex ? 1'h0 : _GEN_14; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_21 = 4'h9 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 105:38 85:27]
  wire  _GEN_22 = 4'h9 == io_BankIndex ? 1'h0 : _GEN_15; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_23 = 4'h9 == io_BankIndex ? 1'h0 : _GEN_16; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_24 = 4'h9 == io_BankIndex ? 1'h0 : _GEN_17; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_25 = 4'h9 == io_BankIndex ? 1'h0 : _GEN_18; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_26 = 4'h9 == io_BankIndex ? 1'h0 : _GEN_19; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_27 = 4'h9 == io_BankIndex ? 1'h0 : _GEN_20; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_28 = 4'h8 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 104:38 84:27]
  wire  _GEN_29 = 4'h8 == io_BankIndex ? 1'h0 : _GEN_21; // @[OuterBuffer.scala 95:24 85:27]
  wire  _GEN_30 = 4'h8 == io_BankIndex ? 1'h0 : _GEN_22; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_31 = 4'h8 == io_BankIndex ? 1'h0 : _GEN_23; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_32 = 4'h8 == io_BankIndex ? 1'h0 : _GEN_24; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_33 = 4'h8 == io_BankIndex ? 1'h0 : _GEN_25; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_34 = 4'h8 == io_BankIndex ? 1'h0 : _GEN_26; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_35 = 4'h8 == io_BankIndex ? 1'h0 : _GEN_27; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_36 = 4'h7 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 103:38 83:27]
  wire  _GEN_37 = 4'h7 == io_BankIndex ? 1'h0 : _GEN_28; // @[OuterBuffer.scala 95:24 84:27]
  wire  _GEN_38 = 4'h7 == io_BankIndex ? 1'h0 : _GEN_29; // @[OuterBuffer.scala 95:24 85:27]
  wire  _GEN_39 = 4'h7 == io_BankIndex ? 1'h0 : _GEN_30; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_40 = 4'h7 == io_BankIndex ? 1'h0 : _GEN_31; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_41 = 4'h7 == io_BankIndex ? 1'h0 : _GEN_32; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_42 = 4'h7 == io_BankIndex ? 1'h0 : _GEN_33; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_43 = 4'h7 == io_BankIndex ? 1'h0 : _GEN_34; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_44 = 4'h7 == io_BankIndex ? 1'h0 : _GEN_35; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_45 = 4'h6 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 102:38 82:27]
  wire  _GEN_46 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_36; // @[OuterBuffer.scala 95:24 83:27]
  wire  _GEN_47 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_37; // @[OuterBuffer.scala 95:24 84:27]
  wire  _GEN_48 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_38; // @[OuterBuffer.scala 95:24 85:27]
  wire  _GEN_49 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_39; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_50 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_40; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_51 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_41; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_52 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_42; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_53 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_43; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_54 = 4'h6 == io_BankIndex ? 1'h0 : _GEN_44; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_55 = 4'h5 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 101:38 81:27]
  wire  _GEN_56 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_45; // @[OuterBuffer.scala 95:24 82:27]
  wire  _GEN_57 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_46; // @[OuterBuffer.scala 95:24 83:27]
  wire  _GEN_58 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_47; // @[OuterBuffer.scala 95:24 84:27]
  wire  _GEN_59 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_48; // @[OuterBuffer.scala 95:24 85:27]
  wire  _GEN_60 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_49; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_61 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_50; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_62 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_51; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_63 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_52; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_64 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_53; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_65 = 4'h5 == io_BankIndex ? 1'h0 : _GEN_54; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_66 = 4'h4 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 100:38 80:27]
  wire  _GEN_67 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_55; // @[OuterBuffer.scala 95:24 81:27]
  wire  _GEN_68 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_56; // @[OuterBuffer.scala 95:24 82:27]
  wire  _GEN_69 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_57; // @[OuterBuffer.scala 95:24 83:27]
  wire  _GEN_70 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_58; // @[OuterBuffer.scala 95:24 84:27]
  wire  _GEN_71 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_59; // @[OuterBuffer.scala 95:24 85:27]
  wire  _GEN_72 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_60; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_73 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_61; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_74 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_62; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_75 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_63; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_76 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_64; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_77 = 4'h4 == io_BankIndex ? 1'h0 : _GEN_65; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_78 = 4'h3 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 79:27 99:38]
  wire  _GEN_79 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_66; // @[OuterBuffer.scala 95:24 80:27]
  wire  _GEN_80 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_67; // @[OuterBuffer.scala 95:24 81:27]
  wire  _GEN_81 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_68; // @[OuterBuffer.scala 95:24 82:27]
  wire  _GEN_82 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_69; // @[OuterBuffer.scala 95:24 83:27]
  wire  _GEN_83 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_70; // @[OuterBuffer.scala 95:24 84:27]
  wire  _GEN_84 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_71; // @[OuterBuffer.scala 95:24 85:27]
  wire  _GEN_85 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_72; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_86 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_73; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_87 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_74; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_88 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_75; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_89 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_76; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_90 = 4'h3 == io_BankIndex ? 1'h0 : _GEN_77; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_91 = 4'h2 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 78:27 98:38]
  wire  _GEN_92 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_78; // @[OuterBuffer.scala 95:24 79:27]
  wire  _GEN_93 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_79; // @[OuterBuffer.scala 95:24 80:27]
  wire  _GEN_94 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_80; // @[OuterBuffer.scala 95:24 81:27]
  wire  _GEN_95 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_81; // @[OuterBuffer.scala 95:24 82:27]
  wire  _GEN_96 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_82; // @[OuterBuffer.scala 95:24 83:27]
  wire  _GEN_97 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_83; // @[OuterBuffer.scala 95:24 84:27]
  wire  _GEN_98 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_84; // @[OuterBuffer.scala 95:24 85:27]
  wire  _GEN_99 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_85; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_100 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_86; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_101 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_87; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_102 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_88; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_103 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_89; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_104 = 4'h2 == io_BankIndex ? 1'h0 : _GEN_90; // @[OuterBuffer.scala 95:24 91:27]
  wire  _GEN_105 = 4'h1 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 77:27 97:38]
  wire  _GEN_106 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_91; // @[OuterBuffer.scala 95:24 78:27]
  wire  _GEN_107 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_92; // @[OuterBuffer.scala 95:24 79:27]
  wire  _GEN_108 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_93; // @[OuterBuffer.scala 95:24 80:27]
  wire  _GEN_109 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_94; // @[OuterBuffer.scala 95:24 81:27]
  wire  _GEN_110 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_95; // @[OuterBuffer.scala 95:24 82:27]
  wire  _GEN_111 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_96; // @[OuterBuffer.scala 95:24 83:27]
  wire  _GEN_112 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_97; // @[OuterBuffer.scala 95:24 84:27]
  wire  _GEN_113 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_98; // @[OuterBuffer.scala 95:24 85:27]
  wire  _GEN_114 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_99; // @[OuterBuffer.scala 95:24 86:27]
  wire  _GEN_115 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_100; // @[OuterBuffer.scala 95:24 87:27]
  wire  _GEN_116 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_101; // @[OuterBuffer.scala 95:24 88:27]
  wire  _GEN_117 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_102; // @[OuterBuffer.scala 95:24 89:27]
  wire  _GEN_118 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_103; // @[OuterBuffer.scala 95:24 90:27]
  wire  _GEN_119 = 4'h1 == io_BankIndex ? 1'h0 : _GEN_104; // @[OuterBuffer.scala 95:24 91:27]
  wire [15:0] _GEN_136 = _T_15 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 131:42 74:27]
  wire [15:0] _GEN_137 = _T_14 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 130:42 73:27]
  wire [15:0] _GEN_138 = _T_14 ? 16'h0 : _GEN_136; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_139 = _T_13 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 129:42 72:27]
  wire [15:0] _GEN_140 = _T_13 ? 16'h0 : _GEN_137; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_141 = _T_13 ? 16'h0 : _GEN_138; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_142 = _T_12 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 128:42 71:27]
  wire [15:0] _GEN_143 = _T_12 ? 16'h0 : _GEN_139; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_144 = _T_12 ? 16'h0 : _GEN_140; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_145 = _T_12 ? 16'h0 : _GEN_141; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_146 = _T_11 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 127:42 70:27]
  wire [15:0] _GEN_147 = _T_11 ? 16'h0 : _GEN_142; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_148 = _T_11 ? 16'h0 : _GEN_143; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_149 = _T_11 ? 16'h0 : _GEN_144; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_150 = _T_11 ? 16'h0 : _GEN_145; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_151 = _T_10 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 126:42 69:27]
  wire [15:0] _GEN_152 = _T_10 ? 16'h0 : _GEN_146; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_153 = _T_10 ? 16'h0 : _GEN_147; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_154 = _T_10 ? 16'h0 : _GEN_148; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_155 = _T_10 ? 16'h0 : _GEN_149; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_156 = _T_10 ? 16'h0 : _GEN_150; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_157 = _T_9 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 125:40 68:27]
  wire [15:0] _GEN_158 = _T_9 ? 16'h0 : _GEN_151; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_159 = _T_9 ? 16'h0 : _GEN_152; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_160 = _T_9 ? 16'h0 : _GEN_153; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_161 = _T_9 ? 16'h0 : _GEN_154; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_162 = _T_9 ? 16'h0 : _GEN_155; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_163 = _T_9 ? 16'h0 : _GEN_156; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_164 = _T_8 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 124:40 67:27]
  wire [15:0] _GEN_165 = _T_8 ? 16'h0 : _GEN_157; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_166 = _T_8 ? 16'h0 : _GEN_158; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_167 = _T_8 ? 16'h0 : _GEN_159; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_168 = _T_8 ? 16'h0 : _GEN_160; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_169 = _T_8 ? 16'h0 : _GEN_161; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_170 = _T_8 ? 16'h0 : _GEN_162; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_171 = _T_8 ? 16'h0 : _GEN_163; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_172 = _T_7 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 123:40 66:27]
  wire [15:0] _GEN_173 = _T_7 ? 16'h0 : _GEN_164; // @[OuterBuffer.scala 115:26 67:27]
  wire [15:0] _GEN_174 = _T_7 ? 16'h0 : _GEN_165; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_175 = _T_7 ? 16'h0 : _GEN_166; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_176 = _T_7 ? 16'h0 : _GEN_167; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_177 = _T_7 ? 16'h0 : _GEN_168; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_178 = _T_7 ? 16'h0 : _GEN_169; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_179 = _T_7 ? 16'h0 : _GEN_170; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_180 = _T_7 ? 16'h0 : _GEN_171; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_181 = _T_6 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 122:40 65:27]
  wire [15:0] _GEN_182 = _T_6 ? 16'h0 : _GEN_172; // @[OuterBuffer.scala 115:26 66:27]
  wire [15:0] _GEN_183 = _T_6 ? 16'h0 : _GEN_173; // @[OuterBuffer.scala 115:26 67:27]
  wire [15:0] _GEN_184 = _T_6 ? 16'h0 : _GEN_174; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_185 = _T_6 ? 16'h0 : _GEN_175; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_186 = _T_6 ? 16'h0 : _GEN_176; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_187 = _T_6 ? 16'h0 : _GEN_177; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_188 = _T_6 ? 16'h0 : _GEN_178; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_189 = _T_6 ? 16'h0 : _GEN_179; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_190 = _T_6 ? 16'h0 : _GEN_180; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_191 = _T_5 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 121:40 64:27]
  wire [15:0] _GEN_192 = _T_5 ? 16'h0 : _GEN_181; // @[OuterBuffer.scala 115:26 65:27]
  wire [15:0] _GEN_193 = _T_5 ? 16'h0 : _GEN_182; // @[OuterBuffer.scala 115:26 66:27]
  wire [15:0] _GEN_194 = _T_5 ? 16'h0 : _GEN_183; // @[OuterBuffer.scala 115:26 67:27]
  wire [15:0] _GEN_195 = _T_5 ? 16'h0 : _GEN_184; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_196 = _T_5 ? 16'h0 : _GEN_185; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_197 = _T_5 ? 16'h0 : _GEN_186; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_198 = _T_5 ? 16'h0 : _GEN_187; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_199 = _T_5 ? 16'h0 : _GEN_188; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_200 = _T_5 ? 16'h0 : _GEN_189; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_201 = _T_5 ? 16'h0 : _GEN_190; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_202 = _T_4 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 120:40 63:27]
  wire [15:0] _GEN_203 = _T_4 ? 16'h0 : _GEN_191; // @[OuterBuffer.scala 115:26 64:27]
  wire [15:0] _GEN_204 = _T_4 ? 16'h0 : _GEN_192; // @[OuterBuffer.scala 115:26 65:27]
  wire [15:0] _GEN_205 = _T_4 ? 16'h0 : _GEN_193; // @[OuterBuffer.scala 115:26 66:27]
  wire [15:0] _GEN_206 = _T_4 ? 16'h0 : _GEN_194; // @[OuterBuffer.scala 115:26 67:27]
  wire [15:0] _GEN_207 = _T_4 ? 16'h0 : _GEN_195; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_208 = _T_4 ? 16'h0 : _GEN_196; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_209 = _T_4 ? 16'h0 : _GEN_197; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_210 = _T_4 ? 16'h0 : _GEN_198; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_211 = _T_4 ? 16'h0 : _GEN_199; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_212 = _T_4 ? 16'h0 : _GEN_200; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_213 = _T_4 ? 16'h0 : _GEN_201; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_214 = _T_3 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 119:40 62:27]
  wire [15:0] _GEN_215 = _T_3 ? 16'h0 : _GEN_202; // @[OuterBuffer.scala 115:26 63:27]
  wire [15:0] _GEN_216 = _T_3 ? 16'h0 : _GEN_203; // @[OuterBuffer.scala 115:26 64:27]
  wire [15:0] _GEN_217 = _T_3 ? 16'h0 : _GEN_204; // @[OuterBuffer.scala 115:26 65:27]
  wire [15:0] _GEN_218 = _T_3 ? 16'h0 : _GEN_205; // @[OuterBuffer.scala 115:26 66:27]
  wire [15:0] _GEN_219 = _T_3 ? 16'h0 : _GEN_206; // @[OuterBuffer.scala 115:26 67:27]
  wire [15:0] _GEN_220 = _T_3 ? 16'h0 : _GEN_207; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_221 = _T_3 ? 16'h0 : _GEN_208; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_222 = _T_3 ? 16'h0 : _GEN_209; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_223 = _T_3 ? 16'h0 : _GEN_210; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_224 = _T_3 ? 16'h0 : _GEN_211; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_225 = _T_3 ? 16'h0 : _GEN_212; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_226 = _T_3 ? 16'h0 : _GEN_213; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_227 = _T_2 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 118:40 61:27]
  wire [15:0] _GEN_228 = _T_2 ? 16'h0 : _GEN_214; // @[OuterBuffer.scala 115:26 62:27]
  wire [15:0] _GEN_229 = _T_2 ? 16'h0 : _GEN_215; // @[OuterBuffer.scala 115:26 63:27]
  wire [15:0] _GEN_230 = _T_2 ? 16'h0 : _GEN_216; // @[OuterBuffer.scala 115:26 64:27]
  wire [15:0] _GEN_231 = _T_2 ? 16'h0 : _GEN_217; // @[OuterBuffer.scala 115:26 65:27]
  wire [15:0] _GEN_232 = _T_2 ? 16'h0 : _GEN_218; // @[OuterBuffer.scala 115:26 66:27]
  wire [15:0] _GEN_233 = _T_2 ? 16'h0 : _GEN_219; // @[OuterBuffer.scala 115:26 67:27]
  wire [15:0] _GEN_234 = _T_2 ? 16'h0 : _GEN_220; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_235 = _T_2 ? 16'h0 : _GEN_221; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_236 = _T_2 ? 16'h0 : _GEN_222; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_237 = _T_2 ? 16'h0 : _GEN_223; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_238 = _T_2 ? 16'h0 : _GEN_224; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_239 = _T_2 ? 16'h0 : _GEN_225; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_240 = _T_2 ? 16'h0 : _GEN_226; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_241 = _T_1 ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 117:40 60:27]
  wire [15:0] _GEN_242 = _T_1 ? 16'h0 : _GEN_227; // @[OuterBuffer.scala 115:26 61:27]
  wire [15:0] _GEN_243 = _T_1 ? 16'h0 : _GEN_228; // @[OuterBuffer.scala 115:26 62:27]
  wire [15:0] _GEN_244 = _T_1 ? 16'h0 : _GEN_229; // @[OuterBuffer.scala 115:26 63:27]
  wire [15:0] _GEN_245 = _T_1 ? 16'h0 : _GEN_230; // @[OuterBuffer.scala 115:26 64:27]
  wire [15:0] _GEN_246 = _T_1 ? 16'h0 : _GEN_231; // @[OuterBuffer.scala 115:26 65:27]
  wire [15:0] _GEN_247 = _T_1 ? 16'h0 : _GEN_232; // @[OuterBuffer.scala 115:26 66:27]
  wire [15:0] _GEN_248 = _T_1 ? 16'h0 : _GEN_233; // @[OuterBuffer.scala 115:26 67:27]
  wire [15:0] _GEN_249 = _T_1 ? 16'h0 : _GEN_234; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_250 = _T_1 ? 16'h0 : _GEN_235; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_251 = _T_1 ? 16'h0 : _GEN_236; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_252 = _T_1 ? 16'h0 : _GEN_237; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_253 = _T_1 ? 16'h0 : _GEN_238; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_254 = _T_1 ? 16'h0 : _GEN_239; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_255 = _T_1 ? 16'h0 : _GEN_240; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_256 = _T ? io_BufferIO_DataIn : 16'h0; // @[OuterBuffer.scala 115:26 116:40 59:27]
  wire [15:0] _GEN_257 = _T ? 16'h0 : _GEN_241; // @[OuterBuffer.scala 115:26 60:27]
  wire [15:0] _GEN_258 = _T ? 16'h0 : _GEN_242; // @[OuterBuffer.scala 115:26 61:27]
  wire [15:0] _GEN_259 = _T ? 16'h0 : _GEN_243; // @[OuterBuffer.scala 115:26 62:27]
  wire [15:0] _GEN_260 = _T ? 16'h0 : _GEN_244; // @[OuterBuffer.scala 115:26 63:27]
  wire [15:0] _GEN_261 = _T ? 16'h0 : _GEN_245; // @[OuterBuffer.scala 115:26 64:27]
  wire [15:0] _GEN_262 = _T ? 16'h0 : _GEN_246; // @[OuterBuffer.scala 115:26 65:27]
  wire [15:0] _GEN_263 = _T ? 16'h0 : _GEN_247; // @[OuterBuffer.scala 115:26 66:27]
  wire [15:0] _GEN_264 = _T ? 16'h0 : _GEN_248; // @[OuterBuffer.scala 115:26 67:27]
  wire [15:0] _GEN_265 = _T ? 16'h0 : _GEN_249; // @[OuterBuffer.scala 115:26 68:27]
  wire [15:0] _GEN_266 = _T ? 16'h0 : _GEN_250; // @[OuterBuffer.scala 115:26 69:27]
  wire [15:0] _GEN_267 = _T ? 16'h0 : _GEN_251; // @[OuterBuffer.scala 115:26 70:27]
  wire [15:0] _GEN_268 = _T ? 16'h0 : _GEN_252; // @[OuterBuffer.scala 115:26 71:27]
  wire [15:0] _GEN_269 = _T ? 16'h0 : _GEN_253; // @[OuterBuffer.scala 115:26 72:27]
  wire [15:0] _GEN_270 = _T ? 16'h0 : _GEN_254; // @[OuterBuffer.scala 115:26 73:27]
  wire [15:0] _GEN_271 = _T ? 16'h0 : _GEN_255; // @[OuterBuffer.scala 115:26 74:27]
  wire [15:0] _GEN_272 = _T_15 ? bank15_io_BankIO_DataOut : 16'h0; // @[OuterBuffer.scala 134:26 150:38 93:23]
  wire [15:0] _GEN_273 = _T_14 ? bank14_io_BankIO_DataOut : _GEN_272; // @[OuterBuffer.scala 134:26 149:38]
  wire [15:0] _GEN_274 = _T_13 ? bank13_io_BankIO_DataOut : _GEN_273; // @[OuterBuffer.scala 134:26 148:38]
  wire [15:0] _GEN_275 = _T_12 ? bank12_io_BankIO_DataOut : _GEN_274; // @[OuterBuffer.scala 134:26 147:38]
  wire [15:0] _GEN_276 = _T_11 ? bank11_io_BankIO_DataOut : _GEN_275; // @[OuterBuffer.scala 134:26 146:38]
  wire [15:0] _GEN_277 = _T_10 ? bank10_io_BankIO_DataOut : _GEN_276; // @[OuterBuffer.scala 134:26 145:38]
  wire [15:0] _GEN_278 = _T_9 ? bank9_io_BankIO_DataOut : _GEN_277; // @[OuterBuffer.scala 134:26 144:37]
  wire [15:0] _GEN_279 = _T_8 ? bank8_io_BankIO_DataOut : _GEN_278; // @[OuterBuffer.scala 134:26 143:37]
  wire [15:0] _GEN_280 = _T_7 ? bank7_io_BankIO_DataOut : _GEN_279; // @[OuterBuffer.scala 134:26 142:37]
  wire [15:0] _GEN_281 = _T_6 ? bank6_io_BankIO_DataOut : _GEN_280; // @[OuterBuffer.scala 134:26 141:37]
  wire [15:0] _GEN_282 = _T_5 ? bank5_io_BankIO_DataOut : _GEN_281; // @[OuterBuffer.scala 134:26 140:37]
  wire [15:0] _GEN_283 = _T_4 ? bank4_io_BankIO_DataOut : _GEN_282; // @[OuterBuffer.scala 134:26 139:37]
  wire [15:0] _GEN_284 = _T_3 ? bank3_io_BankIO_DataOut : _GEN_283; // @[OuterBuffer.scala 134:26 138:37]
  wire [15:0] _GEN_285 = _T_2 ? bank2_io_BankIO_DataOut : _GEN_284; // @[OuterBuffer.scala 134:26 137:37]
  wire [15:0] _GEN_286 = _T_1 ? bank1_io_BankIO_DataOut : _GEN_285; // @[OuterBuffer.scala 134:26 136:37]
  wire [15:0] _GEN_287 = _T ? bank0_io_BankIO_DataOut : _GEN_286; // @[OuterBuffer.scala 134:26 135:37]
  Bank bank0 ( // @[OuterBuffer.scala 41:23]
    .clock(bank0_clock),
    .reset(bank0_reset),
    .io_BankIO_DataIn(bank0_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank0_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank0_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank0_io_BankIO_Enable),
    .io_BankIO_DataOut(bank0_io_BankIO_DataOut)
  );
  Bank bank1 ( // @[OuterBuffer.scala 42:23]
    .clock(bank1_clock),
    .reset(bank1_reset),
    .io_BankIO_DataIn(bank1_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank1_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank1_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank1_io_BankIO_Enable),
    .io_BankIO_DataOut(bank1_io_BankIO_DataOut)
  );
  Bank bank2 ( // @[OuterBuffer.scala 43:23]
    .clock(bank2_clock),
    .reset(bank2_reset),
    .io_BankIO_DataIn(bank2_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank2_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank2_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank2_io_BankIO_Enable),
    .io_BankIO_DataOut(bank2_io_BankIO_DataOut)
  );
  Bank bank3 ( // @[OuterBuffer.scala 44:23]
    .clock(bank3_clock),
    .reset(bank3_reset),
    .io_BankIO_DataIn(bank3_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank3_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank3_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank3_io_BankIO_Enable),
    .io_BankIO_DataOut(bank3_io_BankIO_DataOut)
  );
  Bank bank4 ( // @[OuterBuffer.scala 45:23]
    .clock(bank4_clock),
    .reset(bank4_reset),
    .io_BankIO_DataIn(bank4_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank4_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank4_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank4_io_BankIO_Enable),
    .io_BankIO_DataOut(bank4_io_BankIO_DataOut)
  );
  Bank bank5 ( // @[OuterBuffer.scala 46:23]
    .clock(bank5_clock),
    .reset(bank5_reset),
    .io_BankIO_DataIn(bank5_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank5_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank5_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank5_io_BankIO_Enable),
    .io_BankIO_DataOut(bank5_io_BankIO_DataOut)
  );
  Bank bank6 ( // @[OuterBuffer.scala 47:23]
    .clock(bank6_clock),
    .reset(bank6_reset),
    .io_BankIO_DataIn(bank6_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank6_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank6_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank6_io_BankIO_Enable),
    .io_BankIO_DataOut(bank6_io_BankIO_DataOut)
  );
  Bank bank7 ( // @[OuterBuffer.scala 48:23]
    .clock(bank7_clock),
    .reset(bank7_reset),
    .io_BankIO_DataIn(bank7_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank7_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank7_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank7_io_BankIO_Enable),
    .io_BankIO_DataOut(bank7_io_BankIO_DataOut)
  );
  Bank bank8 ( // @[OuterBuffer.scala 49:23]
    .clock(bank8_clock),
    .reset(bank8_reset),
    .io_BankIO_DataIn(bank8_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank8_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank8_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank8_io_BankIO_Enable),
    .io_BankIO_DataOut(bank8_io_BankIO_DataOut)
  );
  Bank bank9 ( // @[OuterBuffer.scala 50:23]
    .clock(bank9_clock),
    .reset(bank9_reset),
    .io_BankIO_DataIn(bank9_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank9_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank9_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank9_io_BankIO_Enable),
    .io_BankIO_DataOut(bank9_io_BankIO_DataOut)
  );
  Bank bank10 ( // @[OuterBuffer.scala 51:23]
    .clock(bank10_clock),
    .reset(bank10_reset),
    .io_BankIO_DataIn(bank10_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank10_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank10_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank10_io_BankIO_Enable),
    .io_BankIO_DataOut(bank10_io_BankIO_DataOut)
  );
  Bank bank11 ( // @[OuterBuffer.scala 52:23]
    .clock(bank11_clock),
    .reset(bank11_reset),
    .io_BankIO_DataIn(bank11_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank11_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank11_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank11_io_BankIO_Enable),
    .io_BankIO_DataOut(bank11_io_BankIO_DataOut)
  );
  Bank bank12 ( // @[OuterBuffer.scala 53:23]
    .clock(bank12_clock),
    .reset(bank12_reset),
    .io_BankIO_DataIn(bank12_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank12_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank12_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank12_io_BankIO_Enable),
    .io_BankIO_DataOut(bank12_io_BankIO_DataOut)
  );
  Bank bank13 ( // @[OuterBuffer.scala 54:23]
    .clock(bank13_clock),
    .reset(bank13_reset),
    .io_BankIO_DataIn(bank13_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank13_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank13_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank13_io_BankIO_Enable),
    .io_BankIO_DataOut(bank13_io_BankIO_DataOut)
  );
  Bank bank14 ( // @[OuterBuffer.scala 55:23]
    .clock(bank14_clock),
    .reset(bank14_reset),
    .io_BankIO_DataIn(bank14_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank14_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank14_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank14_io_BankIO_Enable),
    .io_BankIO_DataOut(bank14_io_BankIO_DataOut)
  );
  Bank bank15 ( // @[OuterBuffer.scala 56:23]
    .clock(bank15_clock),
    .reset(bank15_reset),
    .io_BankIO_DataIn(bank15_io_BankIO_DataIn),
    .io_BankIO_DataAddr(bank15_io_BankIO_DataAddr),
    .io_BankIO_ReadWrite(bank15_io_BankIO_ReadWrite),
    .io_BankIO_Enable(bank15_io_BankIO_Enable),
    .io_BankIO_DataOut(bank15_io_BankIO_DataOut)
  );
  assign io_BufferIO_DataOut = ~io_BufferIO_ReadWrite ? 16'h0 : _GEN_287; // @[OuterBuffer.scala 114:43 93:23]
  assign bank0_clock = clock;
  assign bank0_reset = reset;
  assign bank0_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_256 : 16'h0; // @[OuterBuffer.scala 114:43 59:27]
  assign bank0_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 154:28]
  assign bank0_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 171:29]
  assign bank0_io_BankIO_Enable = 4'h0 == io_BankIndex & io_BufferIO_Enable; // @[OuterBuffer.scala 95:24 76:27 96:38]
  assign bank1_clock = clock;
  assign bank1_reset = reset;
  assign bank1_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_257 : 16'h0; // @[OuterBuffer.scala 114:43 60:27]
  assign bank1_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 155:28]
  assign bank1_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 172:29]
  assign bank1_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_105; // @[OuterBuffer.scala 95:24 77:27]
  assign bank2_clock = clock;
  assign bank2_reset = reset;
  assign bank2_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_258 : 16'h0; // @[OuterBuffer.scala 114:43 61:27]
  assign bank2_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 156:28]
  assign bank2_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 173:29]
  assign bank2_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_106; // @[OuterBuffer.scala 95:24 78:27]
  assign bank3_clock = clock;
  assign bank3_reset = reset;
  assign bank3_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_259 : 16'h0; // @[OuterBuffer.scala 114:43 62:27]
  assign bank3_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 157:28]
  assign bank3_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 174:29]
  assign bank3_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_107; // @[OuterBuffer.scala 95:24 79:27]
  assign bank4_clock = clock;
  assign bank4_reset = reset;
  assign bank4_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_260 : 16'h0; // @[OuterBuffer.scala 114:43 63:27]
  assign bank4_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 158:28]
  assign bank4_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 175:29]
  assign bank4_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_108; // @[OuterBuffer.scala 95:24 80:27]
  assign bank5_clock = clock;
  assign bank5_reset = reset;
  assign bank5_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_261 : 16'h0; // @[OuterBuffer.scala 114:43 64:27]
  assign bank5_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 159:28]
  assign bank5_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 176:29]
  assign bank5_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_109; // @[OuterBuffer.scala 95:24 81:27]
  assign bank6_clock = clock;
  assign bank6_reset = reset;
  assign bank6_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_262 : 16'h0; // @[OuterBuffer.scala 114:43 65:27]
  assign bank6_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 160:28]
  assign bank6_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 177:29]
  assign bank6_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_110; // @[OuterBuffer.scala 95:24 82:27]
  assign bank7_clock = clock;
  assign bank7_reset = reset;
  assign bank7_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_263 : 16'h0; // @[OuterBuffer.scala 114:43 66:27]
  assign bank7_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 161:28]
  assign bank7_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 178:29]
  assign bank7_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_111; // @[OuterBuffer.scala 95:24 83:27]
  assign bank8_clock = clock;
  assign bank8_reset = reset;
  assign bank8_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_264 : 16'h0; // @[OuterBuffer.scala 114:43 67:27]
  assign bank8_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 162:28]
  assign bank8_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 179:29]
  assign bank8_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_112; // @[OuterBuffer.scala 95:24 84:27]
  assign bank9_clock = clock;
  assign bank9_reset = reset;
  assign bank9_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_265 : 16'h0; // @[OuterBuffer.scala 114:43 68:27]
  assign bank9_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 163:28]
  assign bank9_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 180:29]
  assign bank9_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_113; // @[OuterBuffer.scala 95:24 85:27]
  assign bank10_clock = clock;
  assign bank10_reset = reset;
  assign bank10_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_266 : 16'h0; // @[OuterBuffer.scala 114:43 69:27]
  assign bank10_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 164:29]
  assign bank10_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 181:30]
  assign bank10_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_114; // @[OuterBuffer.scala 95:24 86:27]
  assign bank11_clock = clock;
  assign bank11_reset = reset;
  assign bank11_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_267 : 16'h0; // @[OuterBuffer.scala 114:43 70:27]
  assign bank11_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 165:29]
  assign bank11_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 182:30]
  assign bank11_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_115; // @[OuterBuffer.scala 95:24 87:27]
  assign bank12_clock = clock;
  assign bank12_reset = reset;
  assign bank12_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_268 : 16'h0; // @[OuterBuffer.scala 114:43 71:27]
  assign bank12_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 166:29]
  assign bank12_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 183:30]
  assign bank12_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_116; // @[OuterBuffer.scala 95:24 88:27]
  assign bank13_clock = clock;
  assign bank13_reset = reset;
  assign bank13_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_269 : 16'h0; // @[OuterBuffer.scala 114:43 72:27]
  assign bank13_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 167:29]
  assign bank13_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 184:30]
  assign bank13_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_117; // @[OuterBuffer.scala 95:24 89:27]
  assign bank14_clock = clock;
  assign bank14_reset = reset;
  assign bank14_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_270 : 16'h0; // @[OuterBuffer.scala 114:43 73:27]
  assign bank14_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 168:29]
  assign bank14_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 185:30]
  assign bank14_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_118; // @[OuterBuffer.scala 95:24 90:27]
  assign bank15_clock = clock;
  assign bank15_reset = reset;
  assign bank15_io_BankIO_DataIn = ~io_BufferIO_ReadWrite ? _GEN_271 : 16'h0; // @[OuterBuffer.scala 114:43 74:27]
  assign bank15_io_BankIO_DataAddr = io_BufferIO_DataAddr; // @[OuterBuffer.scala 169:29]
  assign bank15_io_BankIO_ReadWrite = io_BufferIO_ReadWrite; // @[OuterBuffer.scala 186:30]
  assign bank15_io_BankIO_Enable = 4'h0 == io_BankIndex ? 1'h0 : _GEN_119; // @[OuterBuffer.scala 95:24 91:27]
endmodule
module KernelBuffer(
  input         clock,
  input         reset,
  input  [15:0] io_BufferIO_DataIn,
  input  [9:0]  io_BufferIO_DataAddr,
  input         io_BufferIO_ReadWrite,
  input         io_BufferIO_Enable,
  output [15:0] io_BufferIO_DataOut,
  input  [3:0]  io_BankIndex
);
  wire  buf__clock; // @[KernelBuffer.scala 12:19]
  wire  buf__reset; // @[KernelBuffer.scala 12:19]
  wire [15:0] buf__io_BufferIO_DataIn; // @[KernelBuffer.scala 12:19]
  wire [9:0] buf__io_BufferIO_DataAddr; // @[KernelBuffer.scala 12:19]
  wire  buf__io_BufferIO_ReadWrite; // @[KernelBuffer.scala 12:19]
  wire  buf__io_BufferIO_Enable; // @[KernelBuffer.scala 12:19]
  wire [15:0] buf__io_BufferIO_DataOut; // @[KernelBuffer.scala 12:19]
  wire [3:0] buf__io_BankIndex; // @[KernelBuffer.scala 12:19]
  OuterBuffer buf_ ( // @[KernelBuffer.scala 12:19]
    .clock(buf__clock),
    .reset(buf__reset),
    .io_BufferIO_DataIn(buf__io_BufferIO_DataIn),
    .io_BufferIO_DataAddr(buf__io_BufferIO_DataAddr),
    .io_BufferIO_ReadWrite(buf__io_BufferIO_ReadWrite),
    .io_BufferIO_Enable(buf__io_BufferIO_Enable),
    .io_BufferIO_DataOut(buf__io_BufferIO_DataOut),
    .io_BankIndex(buf__io_BankIndex)
  );
  assign io_BufferIO_DataOut = buf__io_BufferIO_DataOut; // @[KernelBuffer.scala 14:15]
  assign buf__clock = clock;
  assign buf__reset = reset;
  assign buf__io_BufferIO_DataIn = io_BufferIO_DataIn; // @[KernelBuffer.scala 14:15]
  assign buf__io_BufferIO_DataAddr = io_BufferIO_DataAddr; // @[KernelBuffer.scala 14:15]
  assign buf__io_BufferIO_ReadWrite = io_BufferIO_ReadWrite; // @[KernelBuffer.scala 14:15]
  assign buf__io_BufferIO_Enable = io_BufferIO_Enable; // @[KernelBuffer.scala 14:15]
  assign buf__io_BankIndex = io_BankIndex; // @[KernelBuffer.scala 15:16]
endmodule
