module AluPool(
  input         clock,
  input         reset,
  input         io_ALUPort_Enable,
  input  [15:0] io_ALUPort_PEDataIn_0,
  input  [15:0] io_ALUPort_PEDataIn_1,
  input  [15:0] io_ALUPort_PEDataIn_2,
  input  [15:0] io_ALUPort_PEDataIn_3,
  input  [15:0] io_ALUPort_PEDataIn_4,
  input  [15:0] io_ALUPort_PEDataIn_5,
  input  [15:0] io_ALUPort_PEDataIn_6,
  input  [15:0] io_ALUPort_PEDataIn_7,
  input  [15:0] io_ALUPort_PEDataIn_8,
  input  [15:0] io_ALUPort_PEDataIn_9,
  input  [15:0] io_ALUPort_PEDataIn_10,
  input  [15:0] io_ALUPort_PEDataIn_11,
  input  [15:0] io_ALUPort_PEDataIn_12,
  input  [15:0] io_ALUPort_PEDataIn_13,
  input  [15:0] io_ALUPort_PEDataIn_14,
  input  [15:0] io_ALUPort_PEDataIn_15,
  output [9:0]  io_ALUPort_Neuron2Addr,
  output [15:0] io_ALUPort_DataOut,
  output [9:0]  io_ALUPort_PsumAddr,
  input  [15:0] io_ALUPort_PsumIn
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] cntMac; // @[AluPool.scala 41:23]
  wire [9:0] _cntMac_T_1 = cntMac + 10'h1; // @[AluPool.scala 45:22]
  wire [16:0] _T_2 = {{1'd0}, io_ALUPort_PEDataIn_0}; // @[AluPool.scala 55:19]
  wire [15:0] _T_5 = _T_2[15:0] + io_ALUPort_PEDataIn_1; // @[AluPool.scala 55:19]
  wire [15:0] _T_7 = _T_5 + io_ALUPort_PEDataIn_2; // @[AluPool.scala 55:19]
  wire [15:0] _T_9 = _T_7 + io_ALUPort_PEDataIn_3; // @[AluPool.scala 55:19]
  wire [15:0] _T_11 = _T_9 + io_ALUPort_PEDataIn_4; // @[AluPool.scala 55:19]
  wire [15:0] _T_13 = _T_11 + io_ALUPort_PEDataIn_5; // @[AluPool.scala 55:19]
  wire [15:0] _T_15 = _T_13 + io_ALUPort_PEDataIn_6; // @[AluPool.scala 55:19]
  wire [15:0] _T_17 = _T_15 + io_ALUPort_PEDataIn_7; // @[AluPool.scala 55:19]
  wire [15:0] _T_19 = _T_17 + io_ALUPort_PEDataIn_8; // @[AluPool.scala 55:19]
  wire [15:0] _T_21 = _T_19 + io_ALUPort_PEDataIn_9; // @[AluPool.scala 55:19]
  wire [15:0] _T_23 = _T_21 + io_ALUPort_PEDataIn_10; // @[AluPool.scala 55:19]
  wire [15:0] _T_25 = _T_23 + io_ALUPort_PEDataIn_11; // @[AluPool.scala 55:19]
  wire [15:0] _T_27 = _T_25 + io_ALUPort_PEDataIn_12; // @[AluPool.scala 55:19]
  wire [15:0] _T_29 = _T_27 + io_ALUPort_PEDataIn_13; // @[AluPool.scala 55:19]
  wire [15:0] _T_31 = _T_29 + io_ALUPort_PEDataIn_14; // @[AluPool.scala 55:19]
  wire [15:0] accumulator = _T_31 + io_ALUPort_PEDataIn_15; // @[AluPool.scala 55:19]
  wire [15:0] _io_ALUPort_DataOut_T_1 = accumulator + io_ALUPort_PsumIn; // @[AluPool.scala 57:39]
  assign io_ALUPort_Neuron2Addr = io_ALUPort_Enable ? cntMac : 10'h0; // @[AluPool.scala 51:38 52:28 59:28]
  assign io_ALUPort_DataOut = io_ALUPort_Enable ? _io_ALUPort_DataOut_T_1 : 16'h0; // @[AluPool.scala 51:38 57:24 61:24]
  assign io_ALUPort_PsumAddr = io_ALUPort_Enable ? cntMac : 10'h0; // @[AluPool.scala 51:38 52:28 59:28]
  always @(posedge clock) begin
    if (reset) begin // @[AluPool.scala 41:23]
      cntMac <= 10'h0; // @[AluPool.scala 41:23]
    end else if (io_ALUPort_Enable) begin // @[AluPool.scala 44:37]
      cntMac <= _cntMac_T_1; // @[AluPool.scala 45:12]
    end else begin
      cntMac <= 10'h0; // @[AluPool.scala 47:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cntMac = _RAND_0[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALUArray(
  input         clock,
  input         reset,
  input         io_ALUPort_0_Enable,
  input  [15:0] io_ALUPort_0_PEDataIn_0,
  input  [15:0] io_ALUPort_0_PEDataIn_1,
  input  [15:0] io_ALUPort_0_PEDataIn_2,
  input  [15:0] io_ALUPort_0_PEDataIn_3,
  input  [15:0] io_ALUPort_0_PEDataIn_4,
  input  [15:0] io_ALUPort_0_PEDataIn_5,
  input  [15:0] io_ALUPort_0_PEDataIn_6,
  input  [15:0] io_ALUPort_0_PEDataIn_7,
  input  [15:0] io_ALUPort_0_PEDataIn_8,
  input  [15:0] io_ALUPort_0_PEDataIn_9,
  input  [15:0] io_ALUPort_0_PEDataIn_10,
  input  [15:0] io_ALUPort_0_PEDataIn_11,
  input  [15:0] io_ALUPort_0_PEDataIn_12,
  input  [15:0] io_ALUPort_0_PEDataIn_13,
  input  [15:0] io_ALUPort_0_PEDataIn_14,
  input  [15:0] io_ALUPort_0_PEDataIn_15,
  output [9:0]  io_ALUPort_0_Neuron2Addr,
  output [3:0]  io_ALUPort_0_BankIdx,
  output [15:0] io_ALUPort_0_DataOut,
  output [9:0]  io_ALUPort_0_PsumAddr,
  input  [15:0] io_ALUPort_0_PsumIn,
  input         io_ALUPort_1_Enable,
  input  [15:0] io_ALUPort_1_PEDataIn_0,
  input  [15:0] io_ALUPort_1_PEDataIn_1,
  input  [15:0] io_ALUPort_1_PEDataIn_2,
  input  [15:0] io_ALUPort_1_PEDataIn_3,
  input  [15:0] io_ALUPort_1_PEDataIn_4,
  input  [15:0] io_ALUPort_1_PEDataIn_5,
  input  [15:0] io_ALUPort_1_PEDataIn_6,
  input  [15:0] io_ALUPort_1_PEDataIn_7,
  input  [15:0] io_ALUPort_1_PEDataIn_8,
  input  [15:0] io_ALUPort_1_PEDataIn_9,
  input  [15:0] io_ALUPort_1_PEDataIn_10,
  input  [15:0] io_ALUPort_1_PEDataIn_11,
  input  [15:0] io_ALUPort_1_PEDataIn_12,
  input  [15:0] io_ALUPort_1_PEDataIn_13,
  input  [15:0] io_ALUPort_1_PEDataIn_14,
  input  [15:0] io_ALUPort_1_PEDataIn_15,
  output [9:0]  io_ALUPort_1_Neuron2Addr,
  output [3:0]  io_ALUPort_1_BankIdx,
  output [15:0] io_ALUPort_1_DataOut,
  output [9:0]  io_ALUPort_1_PsumAddr,
  input  [15:0] io_ALUPort_1_PsumIn,
  input         io_ALUPort_2_Enable,
  input  [15:0] io_ALUPort_2_PEDataIn_0,
  input  [15:0] io_ALUPort_2_PEDataIn_1,
  input  [15:0] io_ALUPort_2_PEDataIn_2,
  input  [15:0] io_ALUPort_2_PEDataIn_3,
  input  [15:0] io_ALUPort_2_PEDataIn_4,
  input  [15:0] io_ALUPort_2_PEDataIn_5,
  input  [15:0] io_ALUPort_2_PEDataIn_6,
  input  [15:0] io_ALUPort_2_PEDataIn_7,
  input  [15:0] io_ALUPort_2_PEDataIn_8,
  input  [15:0] io_ALUPort_2_PEDataIn_9,
  input  [15:0] io_ALUPort_2_PEDataIn_10,
  input  [15:0] io_ALUPort_2_PEDataIn_11,
  input  [15:0] io_ALUPort_2_PEDataIn_12,
  input  [15:0] io_ALUPort_2_PEDataIn_13,
  input  [15:0] io_ALUPort_2_PEDataIn_14,
  input  [15:0] io_ALUPort_2_PEDataIn_15,
  output [9:0]  io_ALUPort_2_Neuron2Addr,
  output [3:0]  io_ALUPort_2_BankIdx,
  output [15:0] io_ALUPort_2_DataOut,
  output [9:0]  io_ALUPort_2_PsumAddr,
  input  [15:0] io_ALUPort_2_PsumIn,
  input         io_ALUPort_3_Enable,
  input  [15:0] io_ALUPort_3_PEDataIn_0,
  input  [15:0] io_ALUPort_3_PEDataIn_1,
  input  [15:0] io_ALUPort_3_PEDataIn_2,
  input  [15:0] io_ALUPort_3_PEDataIn_3,
  input  [15:0] io_ALUPort_3_PEDataIn_4,
  input  [15:0] io_ALUPort_3_PEDataIn_5,
  input  [15:0] io_ALUPort_3_PEDataIn_6,
  input  [15:0] io_ALUPort_3_PEDataIn_7,
  input  [15:0] io_ALUPort_3_PEDataIn_8,
  input  [15:0] io_ALUPort_3_PEDataIn_9,
  input  [15:0] io_ALUPort_3_PEDataIn_10,
  input  [15:0] io_ALUPort_3_PEDataIn_11,
  input  [15:0] io_ALUPort_3_PEDataIn_12,
  input  [15:0] io_ALUPort_3_PEDataIn_13,
  input  [15:0] io_ALUPort_3_PEDataIn_14,
  input  [15:0] io_ALUPort_3_PEDataIn_15,
  output [9:0]  io_ALUPort_3_Neuron2Addr,
  output [3:0]  io_ALUPort_3_BankIdx,
  output [15:0] io_ALUPort_3_DataOut,
  output [9:0]  io_ALUPort_3_PsumAddr,
  input  [15:0] io_ALUPort_3_PsumIn,
  input         io_ALUPort_4_Enable,
  input  [15:0] io_ALUPort_4_PEDataIn_0,
  input  [15:0] io_ALUPort_4_PEDataIn_1,
  input  [15:0] io_ALUPort_4_PEDataIn_2,
  input  [15:0] io_ALUPort_4_PEDataIn_3,
  input  [15:0] io_ALUPort_4_PEDataIn_4,
  input  [15:0] io_ALUPort_4_PEDataIn_5,
  input  [15:0] io_ALUPort_4_PEDataIn_6,
  input  [15:0] io_ALUPort_4_PEDataIn_7,
  input  [15:0] io_ALUPort_4_PEDataIn_8,
  input  [15:0] io_ALUPort_4_PEDataIn_9,
  input  [15:0] io_ALUPort_4_PEDataIn_10,
  input  [15:0] io_ALUPort_4_PEDataIn_11,
  input  [15:0] io_ALUPort_4_PEDataIn_12,
  input  [15:0] io_ALUPort_4_PEDataIn_13,
  input  [15:0] io_ALUPort_4_PEDataIn_14,
  input  [15:0] io_ALUPort_4_PEDataIn_15,
  output [9:0]  io_ALUPort_4_Neuron2Addr,
  output [3:0]  io_ALUPort_4_BankIdx,
  output [15:0] io_ALUPort_4_DataOut,
  output [9:0]  io_ALUPort_4_PsumAddr,
  input  [15:0] io_ALUPort_4_PsumIn,
  input         io_ALUPort_5_Enable,
  input  [15:0] io_ALUPort_5_PEDataIn_0,
  input  [15:0] io_ALUPort_5_PEDataIn_1,
  input  [15:0] io_ALUPort_5_PEDataIn_2,
  input  [15:0] io_ALUPort_5_PEDataIn_3,
  input  [15:0] io_ALUPort_5_PEDataIn_4,
  input  [15:0] io_ALUPort_5_PEDataIn_5,
  input  [15:0] io_ALUPort_5_PEDataIn_6,
  input  [15:0] io_ALUPort_5_PEDataIn_7,
  input  [15:0] io_ALUPort_5_PEDataIn_8,
  input  [15:0] io_ALUPort_5_PEDataIn_9,
  input  [15:0] io_ALUPort_5_PEDataIn_10,
  input  [15:0] io_ALUPort_5_PEDataIn_11,
  input  [15:0] io_ALUPort_5_PEDataIn_12,
  input  [15:0] io_ALUPort_5_PEDataIn_13,
  input  [15:0] io_ALUPort_5_PEDataIn_14,
  input  [15:0] io_ALUPort_5_PEDataIn_15,
  output [9:0]  io_ALUPort_5_Neuron2Addr,
  output [3:0]  io_ALUPort_5_BankIdx,
  output [15:0] io_ALUPort_5_DataOut,
  output [9:0]  io_ALUPort_5_PsumAddr,
  input  [15:0] io_ALUPort_5_PsumIn,
  input         io_ALUPort_6_Enable,
  input  [15:0] io_ALUPort_6_PEDataIn_0,
  input  [15:0] io_ALUPort_6_PEDataIn_1,
  input  [15:0] io_ALUPort_6_PEDataIn_2,
  input  [15:0] io_ALUPort_6_PEDataIn_3,
  input  [15:0] io_ALUPort_6_PEDataIn_4,
  input  [15:0] io_ALUPort_6_PEDataIn_5,
  input  [15:0] io_ALUPort_6_PEDataIn_6,
  input  [15:0] io_ALUPort_6_PEDataIn_7,
  input  [15:0] io_ALUPort_6_PEDataIn_8,
  input  [15:0] io_ALUPort_6_PEDataIn_9,
  input  [15:0] io_ALUPort_6_PEDataIn_10,
  input  [15:0] io_ALUPort_6_PEDataIn_11,
  input  [15:0] io_ALUPort_6_PEDataIn_12,
  input  [15:0] io_ALUPort_6_PEDataIn_13,
  input  [15:0] io_ALUPort_6_PEDataIn_14,
  input  [15:0] io_ALUPort_6_PEDataIn_15,
  output [9:0]  io_ALUPort_6_Neuron2Addr,
  output [3:0]  io_ALUPort_6_BankIdx,
  output [15:0] io_ALUPort_6_DataOut,
  output [9:0]  io_ALUPort_6_PsumAddr,
  input  [15:0] io_ALUPort_6_PsumIn,
  input         io_ALUPort_7_Enable,
  input  [15:0] io_ALUPort_7_PEDataIn_0,
  input  [15:0] io_ALUPort_7_PEDataIn_1,
  input  [15:0] io_ALUPort_7_PEDataIn_2,
  input  [15:0] io_ALUPort_7_PEDataIn_3,
  input  [15:0] io_ALUPort_7_PEDataIn_4,
  input  [15:0] io_ALUPort_7_PEDataIn_5,
  input  [15:0] io_ALUPort_7_PEDataIn_6,
  input  [15:0] io_ALUPort_7_PEDataIn_7,
  input  [15:0] io_ALUPort_7_PEDataIn_8,
  input  [15:0] io_ALUPort_7_PEDataIn_9,
  input  [15:0] io_ALUPort_7_PEDataIn_10,
  input  [15:0] io_ALUPort_7_PEDataIn_11,
  input  [15:0] io_ALUPort_7_PEDataIn_12,
  input  [15:0] io_ALUPort_7_PEDataIn_13,
  input  [15:0] io_ALUPort_7_PEDataIn_14,
  input  [15:0] io_ALUPort_7_PEDataIn_15,
  output [9:0]  io_ALUPort_7_Neuron2Addr,
  output [3:0]  io_ALUPort_7_BankIdx,
  output [15:0] io_ALUPort_7_DataOut,
  output [9:0]  io_ALUPort_7_PsumAddr,
  input  [15:0] io_ALUPort_7_PsumIn,
  input         io_ALUPort_8_Enable,
  input  [15:0] io_ALUPort_8_PEDataIn_0,
  input  [15:0] io_ALUPort_8_PEDataIn_1,
  input  [15:0] io_ALUPort_8_PEDataIn_2,
  input  [15:0] io_ALUPort_8_PEDataIn_3,
  input  [15:0] io_ALUPort_8_PEDataIn_4,
  input  [15:0] io_ALUPort_8_PEDataIn_5,
  input  [15:0] io_ALUPort_8_PEDataIn_6,
  input  [15:0] io_ALUPort_8_PEDataIn_7,
  input  [15:0] io_ALUPort_8_PEDataIn_8,
  input  [15:0] io_ALUPort_8_PEDataIn_9,
  input  [15:0] io_ALUPort_8_PEDataIn_10,
  input  [15:0] io_ALUPort_8_PEDataIn_11,
  input  [15:0] io_ALUPort_8_PEDataIn_12,
  input  [15:0] io_ALUPort_8_PEDataIn_13,
  input  [15:0] io_ALUPort_8_PEDataIn_14,
  input  [15:0] io_ALUPort_8_PEDataIn_15,
  output [9:0]  io_ALUPort_8_Neuron2Addr,
  output [3:0]  io_ALUPort_8_BankIdx,
  output [15:0] io_ALUPort_8_DataOut,
  output [9:0]  io_ALUPort_8_PsumAddr,
  input  [15:0] io_ALUPort_8_PsumIn,
  input         io_ALUPort_9_Enable,
  input  [15:0] io_ALUPort_9_PEDataIn_0,
  input  [15:0] io_ALUPort_9_PEDataIn_1,
  input  [15:0] io_ALUPort_9_PEDataIn_2,
  input  [15:0] io_ALUPort_9_PEDataIn_3,
  input  [15:0] io_ALUPort_9_PEDataIn_4,
  input  [15:0] io_ALUPort_9_PEDataIn_5,
  input  [15:0] io_ALUPort_9_PEDataIn_6,
  input  [15:0] io_ALUPort_9_PEDataIn_7,
  input  [15:0] io_ALUPort_9_PEDataIn_8,
  input  [15:0] io_ALUPort_9_PEDataIn_9,
  input  [15:0] io_ALUPort_9_PEDataIn_10,
  input  [15:0] io_ALUPort_9_PEDataIn_11,
  input  [15:0] io_ALUPort_9_PEDataIn_12,
  input  [15:0] io_ALUPort_9_PEDataIn_13,
  input  [15:0] io_ALUPort_9_PEDataIn_14,
  input  [15:0] io_ALUPort_9_PEDataIn_15,
  output [9:0]  io_ALUPort_9_Neuron2Addr,
  output [3:0]  io_ALUPort_9_BankIdx,
  output [15:0] io_ALUPort_9_DataOut,
  output [9:0]  io_ALUPort_9_PsumAddr,
  input  [15:0] io_ALUPort_9_PsumIn,
  input         io_ALUPort_10_Enable,
  input  [15:0] io_ALUPort_10_PEDataIn_0,
  input  [15:0] io_ALUPort_10_PEDataIn_1,
  input  [15:0] io_ALUPort_10_PEDataIn_2,
  input  [15:0] io_ALUPort_10_PEDataIn_3,
  input  [15:0] io_ALUPort_10_PEDataIn_4,
  input  [15:0] io_ALUPort_10_PEDataIn_5,
  input  [15:0] io_ALUPort_10_PEDataIn_6,
  input  [15:0] io_ALUPort_10_PEDataIn_7,
  input  [15:0] io_ALUPort_10_PEDataIn_8,
  input  [15:0] io_ALUPort_10_PEDataIn_9,
  input  [15:0] io_ALUPort_10_PEDataIn_10,
  input  [15:0] io_ALUPort_10_PEDataIn_11,
  input  [15:0] io_ALUPort_10_PEDataIn_12,
  input  [15:0] io_ALUPort_10_PEDataIn_13,
  input  [15:0] io_ALUPort_10_PEDataIn_14,
  input  [15:0] io_ALUPort_10_PEDataIn_15,
  output [9:0]  io_ALUPort_10_Neuron2Addr,
  output [3:0]  io_ALUPort_10_BankIdx,
  output [15:0] io_ALUPort_10_DataOut,
  output [9:0]  io_ALUPort_10_PsumAddr,
  input  [15:0] io_ALUPort_10_PsumIn,
  input         io_ALUPort_11_Enable,
  input  [15:0] io_ALUPort_11_PEDataIn_0,
  input  [15:0] io_ALUPort_11_PEDataIn_1,
  input  [15:0] io_ALUPort_11_PEDataIn_2,
  input  [15:0] io_ALUPort_11_PEDataIn_3,
  input  [15:0] io_ALUPort_11_PEDataIn_4,
  input  [15:0] io_ALUPort_11_PEDataIn_5,
  input  [15:0] io_ALUPort_11_PEDataIn_6,
  input  [15:0] io_ALUPort_11_PEDataIn_7,
  input  [15:0] io_ALUPort_11_PEDataIn_8,
  input  [15:0] io_ALUPort_11_PEDataIn_9,
  input  [15:0] io_ALUPort_11_PEDataIn_10,
  input  [15:0] io_ALUPort_11_PEDataIn_11,
  input  [15:0] io_ALUPort_11_PEDataIn_12,
  input  [15:0] io_ALUPort_11_PEDataIn_13,
  input  [15:0] io_ALUPort_11_PEDataIn_14,
  input  [15:0] io_ALUPort_11_PEDataIn_15,
  output [9:0]  io_ALUPort_11_Neuron2Addr,
  output [3:0]  io_ALUPort_11_BankIdx,
  output [15:0] io_ALUPort_11_DataOut,
  output [9:0]  io_ALUPort_11_PsumAddr,
  input  [15:0] io_ALUPort_11_PsumIn,
  input         io_ALUPort_12_Enable,
  input  [15:0] io_ALUPort_12_PEDataIn_0,
  input  [15:0] io_ALUPort_12_PEDataIn_1,
  input  [15:0] io_ALUPort_12_PEDataIn_2,
  input  [15:0] io_ALUPort_12_PEDataIn_3,
  input  [15:0] io_ALUPort_12_PEDataIn_4,
  input  [15:0] io_ALUPort_12_PEDataIn_5,
  input  [15:0] io_ALUPort_12_PEDataIn_6,
  input  [15:0] io_ALUPort_12_PEDataIn_7,
  input  [15:0] io_ALUPort_12_PEDataIn_8,
  input  [15:0] io_ALUPort_12_PEDataIn_9,
  input  [15:0] io_ALUPort_12_PEDataIn_10,
  input  [15:0] io_ALUPort_12_PEDataIn_11,
  input  [15:0] io_ALUPort_12_PEDataIn_12,
  input  [15:0] io_ALUPort_12_PEDataIn_13,
  input  [15:0] io_ALUPort_12_PEDataIn_14,
  input  [15:0] io_ALUPort_12_PEDataIn_15,
  output [9:0]  io_ALUPort_12_Neuron2Addr,
  output [3:0]  io_ALUPort_12_BankIdx,
  output [15:0] io_ALUPort_12_DataOut,
  output [9:0]  io_ALUPort_12_PsumAddr,
  input  [15:0] io_ALUPort_12_PsumIn,
  input         io_ALUPort_13_Enable,
  input  [15:0] io_ALUPort_13_PEDataIn_0,
  input  [15:0] io_ALUPort_13_PEDataIn_1,
  input  [15:0] io_ALUPort_13_PEDataIn_2,
  input  [15:0] io_ALUPort_13_PEDataIn_3,
  input  [15:0] io_ALUPort_13_PEDataIn_4,
  input  [15:0] io_ALUPort_13_PEDataIn_5,
  input  [15:0] io_ALUPort_13_PEDataIn_6,
  input  [15:0] io_ALUPort_13_PEDataIn_7,
  input  [15:0] io_ALUPort_13_PEDataIn_8,
  input  [15:0] io_ALUPort_13_PEDataIn_9,
  input  [15:0] io_ALUPort_13_PEDataIn_10,
  input  [15:0] io_ALUPort_13_PEDataIn_11,
  input  [15:0] io_ALUPort_13_PEDataIn_12,
  input  [15:0] io_ALUPort_13_PEDataIn_13,
  input  [15:0] io_ALUPort_13_PEDataIn_14,
  input  [15:0] io_ALUPort_13_PEDataIn_15,
  output [9:0]  io_ALUPort_13_Neuron2Addr,
  output [3:0]  io_ALUPort_13_BankIdx,
  output [15:0] io_ALUPort_13_DataOut,
  output [9:0]  io_ALUPort_13_PsumAddr,
  input  [15:0] io_ALUPort_13_PsumIn,
  input         io_ALUPort_14_Enable,
  input  [15:0] io_ALUPort_14_PEDataIn_0,
  input  [15:0] io_ALUPort_14_PEDataIn_1,
  input  [15:0] io_ALUPort_14_PEDataIn_2,
  input  [15:0] io_ALUPort_14_PEDataIn_3,
  input  [15:0] io_ALUPort_14_PEDataIn_4,
  input  [15:0] io_ALUPort_14_PEDataIn_5,
  input  [15:0] io_ALUPort_14_PEDataIn_6,
  input  [15:0] io_ALUPort_14_PEDataIn_7,
  input  [15:0] io_ALUPort_14_PEDataIn_8,
  input  [15:0] io_ALUPort_14_PEDataIn_9,
  input  [15:0] io_ALUPort_14_PEDataIn_10,
  input  [15:0] io_ALUPort_14_PEDataIn_11,
  input  [15:0] io_ALUPort_14_PEDataIn_12,
  input  [15:0] io_ALUPort_14_PEDataIn_13,
  input  [15:0] io_ALUPort_14_PEDataIn_14,
  input  [15:0] io_ALUPort_14_PEDataIn_15,
  output [9:0]  io_ALUPort_14_Neuron2Addr,
  output [3:0]  io_ALUPort_14_BankIdx,
  output [15:0] io_ALUPort_14_DataOut,
  output [9:0]  io_ALUPort_14_PsumAddr,
  input  [15:0] io_ALUPort_14_PsumIn,
  input         io_ALUPort_15_Enable,
  input  [15:0] io_ALUPort_15_PEDataIn_0,
  input  [15:0] io_ALUPort_15_PEDataIn_1,
  input  [15:0] io_ALUPort_15_PEDataIn_2,
  input  [15:0] io_ALUPort_15_PEDataIn_3,
  input  [15:0] io_ALUPort_15_PEDataIn_4,
  input  [15:0] io_ALUPort_15_PEDataIn_5,
  input  [15:0] io_ALUPort_15_PEDataIn_6,
  input  [15:0] io_ALUPort_15_PEDataIn_7,
  input  [15:0] io_ALUPort_15_PEDataIn_8,
  input  [15:0] io_ALUPort_15_PEDataIn_9,
  input  [15:0] io_ALUPort_15_PEDataIn_10,
  input  [15:0] io_ALUPort_15_PEDataIn_11,
  input  [15:0] io_ALUPort_15_PEDataIn_12,
  input  [15:0] io_ALUPort_15_PEDataIn_13,
  input  [15:0] io_ALUPort_15_PEDataIn_14,
  input  [15:0] io_ALUPort_15_PEDataIn_15,
  output [9:0]  io_ALUPort_15_Neuron2Addr,
  output [3:0]  io_ALUPort_15_BankIdx,
  output [15:0] io_ALUPort_15_DataOut,
  output [9:0]  io_ALUPort_15_PsumAddr,
  input  [15:0] io_ALUPort_15_PsumIn
);
  wire  AluPool_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_1_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_1_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_1_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_1_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_1_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_1_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_2_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_2_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_2_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_2_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_2_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_2_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_3_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_3_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_3_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_3_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_3_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_3_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_4_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_4_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_4_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_4_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_4_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_4_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_5_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_5_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_5_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_5_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_5_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_5_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_6_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_6_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_6_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_6_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_6_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_6_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_7_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_7_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_7_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_7_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_7_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_7_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_8_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_8_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_8_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_8_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_8_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_8_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_9_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_9_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_9_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_9_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_9_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_9_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_10_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_10_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_10_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_10_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_10_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_10_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_11_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_11_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_11_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_11_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_11_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_11_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_12_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_12_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_12_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_12_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_12_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_12_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_13_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_13_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_13_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_13_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_13_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_13_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_14_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_14_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_14_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_14_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_14_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_14_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  wire  AluPool_15_clock; // @[ALUArray.scala 17:51]
  wire  AluPool_15_reset; // @[ALUArray.scala 17:51]
  wire  AluPool_15_io_ALUPort_Enable; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_0; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_1; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_2; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_3; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_4; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_5; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_6; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_7; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_8; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_9; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_10; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_11; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_12; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_13; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_14; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PEDataIn_15; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_15_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_DataOut; // @[ALUArray.scala 17:51]
  wire [9:0] AluPool_15_io_ALUPort_PsumAddr; // @[ALUArray.scala 17:51]
  wire [15:0] AluPool_15_io_ALUPort_PsumIn; // @[ALUArray.scala 17:51]
  AluPool AluPool ( // @[ALUArray.scala 17:51]
    .clock(AluPool_clock),
    .reset(AluPool_reset),
    .io_ALUPort_Enable(AluPool_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_io_ALUPort_PsumIn)
  );
  AluPool AluPool_1 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_1_clock),
    .reset(AluPool_1_reset),
    .io_ALUPort_Enable(AluPool_1_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_1_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_1_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_1_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_1_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_1_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_1_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_1_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_1_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_1_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_1_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_1_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_1_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_1_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_1_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_1_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_1_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_1_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_1_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_1_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_1_io_ALUPort_PsumIn)
  );
  AluPool AluPool_2 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_2_clock),
    .reset(AluPool_2_reset),
    .io_ALUPort_Enable(AluPool_2_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_2_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_2_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_2_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_2_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_2_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_2_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_2_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_2_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_2_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_2_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_2_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_2_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_2_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_2_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_2_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_2_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_2_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_2_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_2_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_2_io_ALUPort_PsumIn)
  );
  AluPool AluPool_3 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_3_clock),
    .reset(AluPool_3_reset),
    .io_ALUPort_Enable(AluPool_3_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_3_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_3_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_3_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_3_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_3_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_3_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_3_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_3_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_3_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_3_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_3_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_3_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_3_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_3_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_3_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_3_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_3_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_3_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_3_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_3_io_ALUPort_PsumIn)
  );
  AluPool AluPool_4 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_4_clock),
    .reset(AluPool_4_reset),
    .io_ALUPort_Enable(AluPool_4_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_4_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_4_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_4_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_4_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_4_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_4_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_4_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_4_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_4_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_4_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_4_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_4_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_4_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_4_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_4_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_4_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_4_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_4_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_4_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_4_io_ALUPort_PsumIn)
  );
  AluPool AluPool_5 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_5_clock),
    .reset(AluPool_5_reset),
    .io_ALUPort_Enable(AluPool_5_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_5_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_5_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_5_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_5_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_5_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_5_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_5_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_5_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_5_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_5_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_5_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_5_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_5_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_5_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_5_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_5_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_5_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_5_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_5_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_5_io_ALUPort_PsumIn)
  );
  AluPool AluPool_6 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_6_clock),
    .reset(AluPool_6_reset),
    .io_ALUPort_Enable(AluPool_6_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_6_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_6_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_6_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_6_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_6_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_6_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_6_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_6_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_6_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_6_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_6_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_6_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_6_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_6_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_6_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_6_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_6_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_6_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_6_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_6_io_ALUPort_PsumIn)
  );
  AluPool AluPool_7 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_7_clock),
    .reset(AluPool_7_reset),
    .io_ALUPort_Enable(AluPool_7_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_7_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_7_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_7_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_7_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_7_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_7_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_7_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_7_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_7_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_7_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_7_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_7_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_7_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_7_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_7_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_7_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_7_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_7_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_7_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_7_io_ALUPort_PsumIn)
  );
  AluPool AluPool_8 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_8_clock),
    .reset(AluPool_8_reset),
    .io_ALUPort_Enable(AluPool_8_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_8_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_8_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_8_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_8_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_8_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_8_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_8_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_8_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_8_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_8_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_8_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_8_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_8_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_8_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_8_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_8_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_8_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_8_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_8_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_8_io_ALUPort_PsumIn)
  );
  AluPool AluPool_9 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_9_clock),
    .reset(AluPool_9_reset),
    .io_ALUPort_Enable(AluPool_9_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_9_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_9_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_9_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_9_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_9_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_9_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_9_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_9_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_9_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_9_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_9_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_9_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_9_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_9_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_9_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_9_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_9_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_9_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_9_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_9_io_ALUPort_PsumIn)
  );
  AluPool AluPool_10 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_10_clock),
    .reset(AluPool_10_reset),
    .io_ALUPort_Enable(AluPool_10_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_10_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_10_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_10_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_10_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_10_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_10_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_10_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_10_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_10_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_10_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_10_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_10_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_10_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_10_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_10_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_10_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_10_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_10_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_10_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_10_io_ALUPort_PsumIn)
  );
  AluPool AluPool_11 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_11_clock),
    .reset(AluPool_11_reset),
    .io_ALUPort_Enable(AluPool_11_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_11_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_11_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_11_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_11_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_11_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_11_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_11_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_11_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_11_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_11_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_11_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_11_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_11_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_11_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_11_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_11_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_11_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_11_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_11_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_11_io_ALUPort_PsumIn)
  );
  AluPool AluPool_12 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_12_clock),
    .reset(AluPool_12_reset),
    .io_ALUPort_Enable(AluPool_12_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_12_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_12_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_12_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_12_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_12_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_12_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_12_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_12_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_12_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_12_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_12_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_12_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_12_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_12_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_12_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_12_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_12_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_12_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_12_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_12_io_ALUPort_PsumIn)
  );
  AluPool AluPool_13 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_13_clock),
    .reset(AluPool_13_reset),
    .io_ALUPort_Enable(AluPool_13_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_13_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_13_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_13_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_13_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_13_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_13_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_13_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_13_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_13_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_13_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_13_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_13_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_13_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_13_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_13_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_13_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_13_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_13_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_13_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_13_io_ALUPort_PsumIn)
  );
  AluPool AluPool_14 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_14_clock),
    .reset(AluPool_14_reset),
    .io_ALUPort_Enable(AluPool_14_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_14_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_14_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_14_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_14_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_14_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_14_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_14_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_14_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_14_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_14_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_14_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_14_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_14_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_14_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_14_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_14_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_14_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_14_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_14_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_14_io_ALUPort_PsumIn)
  );
  AluPool AluPool_15 ( // @[ALUArray.scala 17:51]
    .clock(AluPool_15_clock),
    .reset(AluPool_15_reset),
    .io_ALUPort_Enable(AluPool_15_io_ALUPort_Enable),
    .io_ALUPort_PEDataIn_0(AluPool_15_io_ALUPort_PEDataIn_0),
    .io_ALUPort_PEDataIn_1(AluPool_15_io_ALUPort_PEDataIn_1),
    .io_ALUPort_PEDataIn_2(AluPool_15_io_ALUPort_PEDataIn_2),
    .io_ALUPort_PEDataIn_3(AluPool_15_io_ALUPort_PEDataIn_3),
    .io_ALUPort_PEDataIn_4(AluPool_15_io_ALUPort_PEDataIn_4),
    .io_ALUPort_PEDataIn_5(AluPool_15_io_ALUPort_PEDataIn_5),
    .io_ALUPort_PEDataIn_6(AluPool_15_io_ALUPort_PEDataIn_6),
    .io_ALUPort_PEDataIn_7(AluPool_15_io_ALUPort_PEDataIn_7),
    .io_ALUPort_PEDataIn_8(AluPool_15_io_ALUPort_PEDataIn_8),
    .io_ALUPort_PEDataIn_9(AluPool_15_io_ALUPort_PEDataIn_9),
    .io_ALUPort_PEDataIn_10(AluPool_15_io_ALUPort_PEDataIn_10),
    .io_ALUPort_PEDataIn_11(AluPool_15_io_ALUPort_PEDataIn_11),
    .io_ALUPort_PEDataIn_12(AluPool_15_io_ALUPort_PEDataIn_12),
    .io_ALUPort_PEDataIn_13(AluPool_15_io_ALUPort_PEDataIn_13),
    .io_ALUPort_PEDataIn_14(AluPool_15_io_ALUPort_PEDataIn_14),
    .io_ALUPort_PEDataIn_15(AluPool_15_io_ALUPort_PEDataIn_15),
    .io_ALUPort_Neuron2Addr(AluPool_15_io_ALUPort_Neuron2Addr),
    .io_ALUPort_DataOut(AluPool_15_io_ALUPort_DataOut),
    .io_ALUPort_PsumAddr(AluPool_15_io_ALUPort_PsumAddr),
    .io_ALUPort_PsumIn(AluPool_15_io_ALUPort_PsumIn)
  );
  assign io_ALUPort_0_Neuron2Addr = AluPool_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_0_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_0_DataOut = AluPool_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_0_PsumAddr = AluPool_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_1_Neuron2Addr = AluPool_1_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_1_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_1_DataOut = AluPool_1_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_1_PsumAddr = AluPool_1_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_2_Neuron2Addr = AluPool_2_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_2_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_2_DataOut = AluPool_2_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_2_PsumAddr = AluPool_2_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_3_Neuron2Addr = AluPool_3_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_3_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_3_DataOut = AluPool_3_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_3_PsumAddr = AluPool_3_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_4_Neuron2Addr = AluPool_4_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_4_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_4_DataOut = AluPool_4_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_4_PsumAddr = AluPool_4_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_5_Neuron2Addr = AluPool_5_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_5_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_5_DataOut = AluPool_5_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_5_PsumAddr = AluPool_5_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_6_Neuron2Addr = AluPool_6_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_6_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_6_DataOut = AluPool_6_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_6_PsumAddr = AluPool_6_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_7_Neuron2Addr = AluPool_7_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_7_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_7_DataOut = AluPool_7_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_7_PsumAddr = AluPool_7_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_8_Neuron2Addr = AluPool_8_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_8_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_8_DataOut = AluPool_8_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_8_PsumAddr = AluPool_8_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_9_Neuron2Addr = AluPool_9_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_9_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_9_DataOut = AluPool_9_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_9_PsumAddr = AluPool_9_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_10_Neuron2Addr = AluPool_10_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_10_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_10_DataOut = AluPool_10_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_10_PsumAddr = AluPool_10_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_11_Neuron2Addr = AluPool_11_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_11_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_11_DataOut = AluPool_11_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_11_PsumAddr = AluPool_11_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_12_Neuron2Addr = AluPool_12_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_12_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_12_DataOut = AluPool_12_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_12_PsumAddr = AluPool_12_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_13_Neuron2Addr = AluPool_13_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_13_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_13_DataOut = AluPool_13_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_13_PsumAddr = AluPool_13_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_14_Neuron2Addr = AluPool_14_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_14_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_14_DataOut = AluPool_14_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_14_PsumAddr = AluPool_14_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_15_Neuron2Addr = AluPool_15_io_ALUPort_Neuron2Addr; // @[ALUArray.scala 24:31]
  assign io_ALUPort_15_BankIdx = 4'h0; // @[ALUArray.scala 24:31]
  assign io_ALUPort_15_DataOut = AluPool_15_io_ALUPort_DataOut; // @[ALUArray.scala 24:31]
  assign io_ALUPort_15_PsumAddr = AluPool_15_io_ALUPort_PsumAddr; // @[ALUArray.scala 24:31]
  assign AluPool_clock = clock;
  assign AluPool_reset = reset;
  assign AluPool_io_ALUPort_Enable = io_ALUPort_0_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_0 = io_ALUPort_0_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_1 = io_ALUPort_0_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_2 = io_ALUPort_0_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_3 = io_ALUPort_0_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_4 = io_ALUPort_0_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_5 = io_ALUPort_0_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_6 = io_ALUPort_0_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_7 = io_ALUPort_0_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_8 = io_ALUPort_0_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_9 = io_ALUPort_0_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_10 = io_ALUPort_0_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_11 = io_ALUPort_0_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_12 = io_ALUPort_0_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_13 = io_ALUPort_0_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_14 = io_ALUPort_0_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PEDataIn_15 = io_ALUPort_0_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_io_ALUPort_PsumIn = io_ALUPort_0_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_1_clock = clock;
  assign AluPool_1_reset = reset;
  assign AluPool_1_io_ALUPort_Enable = io_ALUPort_1_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_0 = io_ALUPort_1_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_1 = io_ALUPort_1_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_2 = io_ALUPort_1_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_3 = io_ALUPort_1_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_4 = io_ALUPort_1_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_5 = io_ALUPort_1_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_6 = io_ALUPort_1_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_7 = io_ALUPort_1_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_8 = io_ALUPort_1_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_9 = io_ALUPort_1_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_10 = io_ALUPort_1_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_11 = io_ALUPort_1_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_12 = io_ALUPort_1_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_13 = io_ALUPort_1_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_14 = io_ALUPort_1_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PEDataIn_15 = io_ALUPort_1_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_1_io_ALUPort_PsumIn = io_ALUPort_1_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_2_clock = clock;
  assign AluPool_2_reset = reset;
  assign AluPool_2_io_ALUPort_Enable = io_ALUPort_2_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_0 = io_ALUPort_2_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_1 = io_ALUPort_2_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_2 = io_ALUPort_2_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_3 = io_ALUPort_2_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_4 = io_ALUPort_2_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_5 = io_ALUPort_2_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_6 = io_ALUPort_2_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_7 = io_ALUPort_2_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_8 = io_ALUPort_2_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_9 = io_ALUPort_2_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_10 = io_ALUPort_2_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_11 = io_ALUPort_2_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_12 = io_ALUPort_2_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_13 = io_ALUPort_2_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_14 = io_ALUPort_2_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PEDataIn_15 = io_ALUPort_2_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_2_io_ALUPort_PsumIn = io_ALUPort_2_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_3_clock = clock;
  assign AluPool_3_reset = reset;
  assign AluPool_3_io_ALUPort_Enable = io_ALUPort_3_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_0 = io_ALUPort_3_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_1 = io_ALUPort_3_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_2 = io_ALUPort_3_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_3 = io_ALUPort_3_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_4 = io_ALUPort_3_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_5 = io_ALUPort_3_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_6 = io_ALUPort_3_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_7 = io_ALUPort_3_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_8 = io_ALUPort_3_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_9 = io_ALUPort_3_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_10 = io_ALUPort_3_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_11 = io_ALUPort_3_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_12 = io_ALUPort_3_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_13 = io_ALUPort_3_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_14 = io_ALUPort_3_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PEDataIn_15 = io_ALUPort_3_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_3_io_ALUPort_PsumIn = io_ALUPort_3_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_4_clock = clock;
  assign AluPool_4_reset = reset;
  assign AluPool_4_io_ALUPort_Enable = io_ALUPort_4_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_0 = io_ALUPort_4_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_1 = io_ALUPort_4_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_2 = io_ALUPort_4_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_3 = io_ALUPort_4_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_4 = io_ALUPort_4_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_5 = io_ALUPort_4_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_6 = io_ALUPort_4_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_7 = io_ALUPort_4_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_8 = io_ALUPort_4_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_9 = io_ALUPort_4_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_10 = io_ALUPort_4_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_11 = io_ALUPort_4_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_12 = io_ALUPort_4_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_13 = io_ALUPort_4_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_14 = io_ALUPort_4_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PEDataIn_15 = io_ALUPort_4_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_4_io_ALUPort_PsumIn = io_ALUPort_4_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_5_clock = clock;
  assign AluPool_5_reset = reset;
  assign AluPool_5_io_ALUPort_Enable = io_ALUPort_5_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_0 = io_ALUPort_5_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_1 = io_ALUPort_5_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_2 = io_ALUPort_5_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_3 = io_ALUPort_5_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_4 = io_ALUPort_5_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_5 = io_ALUPort_5_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_6 = io_ALUPort_5_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_7 = io_ALUPort_5_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_8 = io_ALUPort_5_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_9 = io_ALUPort_5_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_10 = io_ALUPort_5_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_11 = io_ALUPort_5_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_12 = io_ALUPort_5_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_13 = io_ALUPort_5_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_14 = io_ALUPort_5_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PEDataIn_15 = io_ALUPort_5_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_5_io_ALUPort_PsumIn = io_ALUPort_5_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_6_clock = clock;
  assign AluPool_6_reset = reset;
  assign AluPool_6_io_ALUPort_Enable = io_ALUPort_6_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_0 = io_ALUPort_6_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_1 = io_ALUPort_6_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_2 = io_ALUPort_6_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_3 = io_ALUPort_6_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_4 = io_ALUPort_6_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_5 = io_ALUPort_6_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_6 = io_ALUPort_6_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_7 = io_ALUPort_6_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_8 = io_ALUPort_6_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_9 = io_ALUPort_6_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_10 = io_ALUPort_6_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_11 = io_ALUPort_6_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_12 = io_ALUPort_6_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_13 = io_ALUPort_6_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_14 = io_ALUPort_6_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PEDataIn_15 = io_ALUPort_6_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_6_io_ALUPort_PsumIn = io_ALUPort_6_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_7_clock = clock;
  assign AluPool_7_reset = reset;
  assign AluPool_7_io_ALUPort_Enable = io_ALUPort_7_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_0 = io_ALUPort_7_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_1 = io_ALUPort_7_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_2 = io_ALUPort_7_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_3 = io_ALUPort_7_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_4 = io_ALUPort_7_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_5 = io_ALUPort_7_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_6 = io_ALUPort_7_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_7 = io_ALUPort_7_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_8 = io_ALUPort_7_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_9 = io_ALUPort_7_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_10 = io_ALUPort_7_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_11 = io_ALUPort_7_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_12 = io_ALUPort_7_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_13 = io_ALUPort_7_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_14 = io_ALUPort_7_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PEDataIn_15 = io_ALUPort_7_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_7_io_ALUPort_PsumIn = io_ALUPort_7_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_8_clock = clock;
  assign AluPool_8_reset = reset;
  assign AluPool_8_io_ALUPort_Enable = io_ALUPort_8_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_0 = io_ALUPort_8_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_1 = io_ALUPort_8_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_2 = io_ALUPort_8_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_3 = io_ALUPort_8_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_4 = io_ALUPort_8_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_5 = io_ALUPort_8_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_6 = io_ALUPort_8_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_7 = io_ALUPort_8_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_8 = io_ALUPort_8_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_9 = io_ALUPort_8_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_10 = io_ALUPort_8_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_11 = io_ALUPort_8_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_12 = io_ALUPort_8_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_13 = io_ALUPort_8_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_14 = io_ALUPort_8_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PEDataIn_15 = io_ALUPort_8_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_8_io_ALUPort_PsumIn = io_ALUPort_8_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_9_clock = clock;
  assign AluPool_9_reset = reset;
  assign AluPool_9_io_ALUPort_Enable = io_ALUPort_9_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_0 = io_ALUPort_9_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_1 = io_ALUPort_9_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_2 = io_ALUPort_9_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_3 = io_ALUPort_9_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_4 = io_ALUPort_9_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_5 = io_ALUPort_9_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_6 = io_ALUPort_9_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_7 = io_ALUPort_9_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_8 = io_ALUPort_9_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_9 = io_ALUPort_9_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_10 = io_ALUPort_9_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_11 = io_ALUPort_9_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_12 = io_ALUPort_9_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_13 = io_ALUPort_9_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_14 = io_ALUPort_9_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PEDataIn_15 = io_ALUPort_9_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_9_io_ALUPort_PsumIn = io_ALUPort_9_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_10_clock = clock;
  assign AluPool_10_reset = reset;
  assign AluPool_10_io_ALUPort_Enable = io_ALUPort_10_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_0 = io_ALUPort_10_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_1 = io_ALUPort_10_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_2 = io_ALUPort_10_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_3 = io_ALUPort_10_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_4 = io_ALUPort_10_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_5 = io_ALUPort_10_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_6 = io_ALUPort_10_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_7 = io_ALUPort_10_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_8 = io_ALUPort_10_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_9 = io_ALUPort_10_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_10 = io_ALUPort_10_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_11 = io_ALUPort_10_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_12 = io_ALUPort_10_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_13 = io_ALUPort_10_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_14 = io_ALUPort_10_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PEDataIn_15 = io_ALUPort_10_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_10_io_ALUPort_PsumIn = io_ALUPort_10_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_11_clock = clock;
  assign AluPool_11_reset = reset;
  assign AluPool_11_io_ALUPort_Enable = io_ALUPort_11_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_0 = io_ALUPort_11_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_1 = io_ALUPort_11_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_2 = io_ALUPort_11_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_3 = io_ALUPort_11_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_4 = io_ALUPort_11_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_5 = io_ALUPort_11_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_6 = io_ALUPort_11_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_7 = io_ALUPort_11_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_8 = io_ALUPort_11_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_9 = io_ALUPort_11_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_10 = io_ALUPort_11_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_11 = io_ALUPort_11_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_12 = io_ALUPort_11_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_13 = io_ALUPort_11_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_14 = io_ALUPort_11_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PEDataIn_15 = io_ALUPort_11_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_11_io_ALUPort_PsumIn = io_ALUPort_11_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_12_clock = clock;
  assign AluPool_12_reset = reset;
  assign AluPool_12_io_ALUPort_Enable = io_ALUPort_12_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_0 = io_ALUPort_12_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_1 = io_ALUPort_12_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_2 = io_ALUPort_12_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_3 = io_ALUPort_12_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_4 = io_ALUPort_12_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_5 = io_ALUPort_12_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_6 = io_ALUPort_12_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_7 = io_ALUPort_12_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_8 = io_ALUPort_12_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_9 = io_ALUPort_12_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_10 = io_ALUPort_12_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_11 = io_ALUPort_12_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_12 = io_ALUPort_12_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_13 = io_ALUPort_12_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_14 = io_ALUPort_12_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PEDataIn_15 = io_ALUPort_12_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_12_io_ALUPort_PsumIn = io_ALUPort_12_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_13_clock = clock;
  assign AluPool_13_reset = reset;
  assign AluPool_13_io_ALUPort_Enable = io_ALUPort_13_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_0 = io_ALUPort_13_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_1 = io_ALUPort_13_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_2 = io_ALUPort_13_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_3 = io_ALUPort_13_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_4 = io_ALUPort_13_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_5 = io_ALUPort_13_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_6 = io_ALUPort_13_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_7 = io_ALUPort_13_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_8 = io_ALUPort_13_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_9 = io_ALUPort_13_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_10 = io_ALUPort_13_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_11 = io_ALUPort_13_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_12 = io_ALUPort_13_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_13 = io_ALUPort_13_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_14 = io_ALUPort_13_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PEDataIn_15 = io_ALUPort_13_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_13_io_ALUPort_PsumIn = io_ALUPort_13_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_14_clock = clock;
  assign AluPool_14_reset = reset;
  assign AluPool_14_io_ALUPort_Enable = io_ALUPort_14_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_0 = io_ALUPort_14_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_1 = io_ALUPort_14_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_2 = io_ALUPort_14_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_3 = io_ALUPort_14_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_4 = io_ALUPort_14_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_5 = io_ALUPort_14_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_6 = io_ALUPort_14_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_7 = io_ALUPort_14_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_8 = io_ALUPort_14_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_9 = io_ALUPort_14_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_10 = io_ALUPort_14_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_11 = io_ALUPort_14_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_12 = io_ALUPort_14_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_13 = io_ALUPort_14_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_14 = io_ALUPort_14_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PEDataIn_15 = io_ALUPort_14_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_14_io_ALUPort_PsumIn = io_ALUPort_14_PsumIn; // @[ALUArray.scala 24:31]
  assign AluPool_15_clock = clock;
  assign AluPool_15_reset = reset;
  assign AluPool_15_io_ALUPort_Enable = io_ALUPort_15_Enable; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_0 = io_ALUPort_15_PEDataIn_0; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_1 = io_ALUPort_15_PEDataIn_1; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_2 = io_ALUPort_15_PEDataIn_2; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_3 = io_ALUPort_15_PEDataIn_3; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_4 = io_ALUPort_15_PEDataIn_4; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_5 = io_ALUPort_15_PEDataIn_5; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_6 = io_ALUPort_15_PEDataIn_6; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_7 = io_ALUPort_15_PEDataIn_7; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_8 = io_ALUPort_15_PEDataIn_8; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_9 = io_ALUPort_15_PEDataIn_9; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_10 = io_ALUPort_15_PEDataIn_10; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_11 = io_ALUPort_15_PEDataIn_11; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_12 = io_ALUPort_15_PEDataIn_12; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_13 = io_ALUPort_15_PEDataIn_13; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_14 = io_ALUPort_15_PEDataIn_14; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PEDataIn_15 = io_ALUPort_15_PEDataIn_15; // @[ALUArray.scala 24:31]
  assign AluPool_15_io_ALUPort_PsumIn = io_ALUPort_15_PsumIn; // @[ALUArray.scala 24:31]
endmodule
